�csklearn.ensemble._forest
RandomForestClassifier
q )�q}q(X   base_estimatorqcsklearn.tree._classes
DecisionTreeClassifier
q)�q}q(X	   criterionqX   giniqX   splitterq	X   bestq
X	   max_depthqNX   min_samples_splitqKX   min_samples_leafqKX   min_weight_fraction_leafqG        X   max_featuresqNX   max_leaf_nodesqNX   random_stateqNX   min_impurity_decreaseqG        X   class_weightqNX	   ccp_alphaqG        X   _sklearn_versionqX   1.0.2qubX   n_estimatorsqKX   estimator_paramsq(hhhhhhhhhhtqX	   bootstrapq�X	   oob_scoreq�X   n_jobsqNhK X   verboseqK X
   warm_startq�hNX   max_samplesqNhhhNhKhKhG        hX   autoq hNhG        hG        X   feature_names_in_q!cnumpy.core.multiarray
_reconstruct
q"cnumpy
ndarray
q#K �q$Cbq%�q&Rq'(KK�q(cnumpy
dtype
q)X   O8q*���q+Rq,(KX   |q-NNNJ����J����K?tq.b�]q/(X   Ageq0X   Sexq1X   ChestPainTypeq2X	   RestingBPq3X   Cholesterolq4X	   FastingBSq5X
   RestingECGq6X   MaxHRq7X   ExerciseAnginaq8X   Oldpeakq9X   ST_Slopeq:etq;bX   n_features_in_q<KX
   n_outputs_q=KX   classes_q>h"h#K �q?h%�q@RqA(KK�qBh)X   i8qC���qDRqE(KX   <qFNNNJ����J����K tqGb�C               qHtqIbX
   n_classes_qJKX   base_estimator_qKhX   estimators_qL]qM(h)�qN}qO(hhh	h
hNhKhKhG        hh hNhJ�
hG        hNhG        h<Kh=Kh>h"h#K �qPh%�qQRqR(KK�qSh)X   f8qT���qURqV(KhFNNNJ����J����K tqWb�C              �?qXtqYbhJcnumpy.core.multiarray
scalar
qZhEC       q[�q\Rq]X   max_features_q^KX   tree_q_csklearn.tree._tree
Tree
q`Kh"h#K �qah%�qbRqc(KK�qdhE�C       qetqfbK�qgRqh}qi(hKX
   node_countqjK�X   nodesqkh"h#K �qlh%�qmRqn(KK��qoh)X   V56qp���qqRqr(Kh-N(X
   left_childqsX   right_childqtX   featurequX	   thresholdqvX   impurityqwX   n_node_samplesqxX   weighted_n_node_samplesqytqz}q{(hsh)X   i8q|���q}Rq~(KhFNNNJ����J����K tqbK �q�hth~K�q�huh~K�q�hvhVK�q�hwhVK �q�hxh~K(�q�hyhVK0�q�uK8KKtq�b�BX7         �                    �?j8je3�?�           ��@       e                    �?�}�	���?           �y@       R                   �a@��k=.��?�            �t@       %                   `a@0`�#��?�             n@               	          ����?p�"�0�?X            �b@                          `_@���^��?9            @X@                          �_@0�й���?*            @R@              
             �?�7��?            �C@	       
                    �?      �?             @������������������������       �                     �?������������������������       �                     @                          xr@��?^�k�?            �A@������������������������       �                     A@������������������������       �                     �?                          �[@H�V�e��?             A@                           �M@p�ݯ��?             3@                          �Z@      �?             ,@                          �V@�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     .@                           @H@�q�q�?             8@������������������������       �                     "@                           �O@��S���?
             .@                            L@�n_Y�K�?	             *@              	             �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @!       "                   �`@ pƵHP�?             J@������������������������       �                     E@#       $                   @M@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@&       =       	          ����? �.�6��?:             W@'       <                   �e@N{�T6�?$            �K@(       ;                    �?(옄��?!             G@)       4                   �_@�K��&�?            �E@*       -                   Pb@��}*_��?             ;@+       ,                   �^@      �?              @������������������������       �                     @������������������������       �                      @.       1                    �?���y4F�?             3@/       0                   �c@      �?             @������������������������       �                     �?������������������������       �                     @2       3                    �B@��S�ۿ?             .@������������������������       �                     �?������������������������       �        
             ,@5       6                   `a@      �?
             0@������������������������       �                     "@7       :                   g@؇���X�?             @8       9                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     "@>       E                   @j@��G���?            �B@?       D                   �h@      �?              @@       C                   �d@�q�q�?             @A       B                    �E@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @F       G                    �?ܷ��?��?             =@������������������������       �                     $@H       M                    �?�S����?             3@I       J                   �c@r�q��?             @������������������������       �                     @K       L       	          033�?      �?              @������������������������       �                     �?������������������������       �                     �?N       O                   0c@8�Z$���?             *@������������������������       �                     $@P       Q                   `n@�q�q�?             @������������������������       �                     �?������������������������       �                      @S       d                    �R@���7�?6             V@T       [                    �H@XB���?5            �U@U       X                    �?�r����?
             .@V       W       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?Y       Z                   �w@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?\       ]       	          033@�k~X��?+             R@������������������������       �                    �G@^       _                   �`@`2U0*��?             9@������������������������       �                     (@`       c                   Pm@$�q-�?             *@a       b                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?f                          �`@U7W1�?9            �T@g       r                    �I@�zv�X�?             F@h       i       	          ������q�q�?             2@������������������������       �                      @j       o                   �b@      �?
             0@k       n                    @E@r�q��?             (@l       m                   �U@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@p       q                    �?      �?             @������������������������       �                      @������������������������       �                      @s       x                    `@���B���?             :@t       w       	          @33�?�t����?
             1@u       v                   @W@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @������������������������       �                      @y       ~                    �?�q�q�?             "@z       }                   �\@      �?             @{       |                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   pb@��-�=��?            �C@������������������������       �                     1@�       �                    �M@"pc�
�?             6@�       �                   �]@���Q��?             $@������������������������       �                     @�       �                   `_@z�G�z�?             @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        	             (@�       �                    @K@"\�����?�             t@�       �                    @��2(&�?x             f@�       �                    �?3��e��?r            �d@�       �                   `l@��	,UP�?=             W@������������������������       �                     B@�       �                   �[@4և����?%             L@�       �                    �I@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   pg@ ��WV�?"             J@�       �                    �?���J��?!            �I@�       �       	          hff @�Ń��̧?             E@������������������������       �                    �D@������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?�       �                    �?�7�QJW�?5            �R@�       �                    T@ ����?0            @P@�       �                    �?���Q��?             @�       �                   �`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �       
             �?��S�ۿ?-             N@������������������������       �                     0@�       �                   @^@�C��2(�?"             F@�       �                    �?�S����?             3@������������������������       �                     @�       �                    @H@      �?
             (@������������������������       �                     @�       �                   �n@և���X�?             @�       �                   @a@�q�q�?             @������������������������       �                      @�       �                     I@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                    b@`2U0*��?             9@�       �                    �H@ףp=
�?             $@������������������������       �                     @�       �                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     .@�       �                    @I@���Q��?             $@������������������������       �                     @������������������������       �                     @�       �                    �?�q�q�?             "@�       �                   pd@���Q��?             @������������������������       �                     �?�       �                    �C@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       
             �?      �?X            @b@�       �                    \@��7	C)�?C            @Z@�       �                    `@r�q��?             2@������������������������       �                     "@�       �                    @�q�q�?             "@�       �                    l@؇���X�?             @�       �                   �U@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �       	          033�?�q�q�?7            �U@�       �                    �?z�G�z�?/            �Q@������������������������       �                     1@�       �                   �q@Ȩ�I��?"            �J@�       �                   �O@�����?            �H@�       �                    �P@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �?(L���?            �E@�       �                   �`@     ��?
             0@�       �                    d@�z�G��?             $@�       �                    �M@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                     P@�����H�?             ;@�       �                    d@ �q�q�?             8@������������������������       �        	             .@�       �                    @�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                    �?�q�q�?             @�       �                   `a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?�t����?             1@������������������������       �                      @������������������������       �                     .@�       �       	          833�?������?            �D@�       �                   Pa@�C��2(�?             &@������������������������       �                     @�       �                    `@r�q��?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?��S�ۿ?             >@�       �                    �?r�q��?             @������������������������       �                      @�       �                   �Y@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �? �q�q�?	             8@������������������������       �                     @�       �       	             @P���Q�?             4@������������������������       �                     3@������������������������       �                     �?q�tq�bX   valuesq�h"h#K �q�h%�q�Rq�(KK�KK�q�hV�B�       Ps@     �z@      U@     �t@     �O@     �p@     �M@     �f@      2@     ``@      1@      T@      "@      P@       @     �B@      �?      @      �?                      @      �?      A@              A@      �?              @      ;@      @      (@      @      @      @      @      @                      @      @                      @              .@       @      0@              "@       @      @       @      @      @      @      @                      @      @                       @      �?     �I@              E@      �?      "@      �?                      "@     �D@     �I@      A@      5@      9@      5@      9@      2@      $@      1@      @       @      @                       @      @      .@      @      �?              �?      @              �?      ,@      �?                      ,@      .@      �?      "@              @      �?      �?      �?      �?                      �?      @                      @      "@              @      >@      @      @       @      @       @      �?              �?       @                      @       @              @      :@              $@      @      0@      �?      @              @      �?      �?      �?                      �?       @      &@              $@       @      �?              �?       @              @      U@      @      U@       @      *@      �?      �?      �?                      �?      �?      (@              (@      �?              �?     �Q@             �G@      �?      8@              (@      �?      (@      �?      @              @      �?                      "@      �?              5@      O@      1@      ;@      (@      @               @      (@      @      $@       @      �?       @      �?                       @      "@               @       @       @                       @      @      5@       @      .@       @      @       @                      @               @      @      @      @      �?      �?      �?      �?                      �?       @                      @      @     �A@              1@      @      2@      @      @              @      @      �?      �?      �?      �?                      �?      @                      (@      l@     @X@      c@      8@     �b@      2@     �U@      @      B@             �I@      @      �?      @              @      �?              I@       @      I@      �?     �D@      �?     �D@                      �?      "@                      �?      O@      *@      M@      @       @      @       @       @       @                       @              �?      L@      @      0@              D@      @      0@      @      @              "@      @      @              @      @      @       @       @               @       @               @       @                      �?      8@      �?      "@      �?      @               @      �?       @                      �?      .@              @      @              @      @              @      @      @       @              �?      @      �?              �?      @                      @     @R@     @R@     �N@      F@      @      .@              "@      @      @      �?      @      �?      �?              �?      �?                      @       @              M@      =@      L@      ,@      1@             �C@      ,@     �C@      $@       @      @              @       @             �B@      @      *@      @      @      @       @      @              @       @              @              @              8@      @      7@      �?      .@               @      �?       @                      �?      �?       @      �?      �?      �?                      �?              �?              @       @      .@       @                      .@      (@      =@      $@      �?      @              @      �?      @              �?      �?      �?                      �?       @      <@      �?      @               @      �?      @      �?                      @      �?      7@              @      �?      3@              3@      �?        q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ/��hG        hNhG        h<Kh=Kh>h"h#K �q�h%�q�Rq�(KK�q�hV�C              �?q�tq�bhJhZhEC       q��q�Rq�h^Kh_h`Kh"h#K �q�h%�q�Rq�(KK�q�hE�C       q�tq�bK�q�Rq�}q�(hKhjK�hkh"h#K �q�h%�q�Rq�(KK��q�hr�Bx6         �       	          ����?4�5����?�           ��@       9                    �?�N2��?�            �w@                          @E@��7�G%�?Y             c@              
             �?�˹�m��?             C@                           �?XB���?             =@                           �H@�C��2(�?             &@������������������������       �                     @       	       
             �?      �?             @������������������������       �                     �?
                          �_@�q�q�?             @������������������������       �                     �?                          �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             2@                           �?�<ݚ�?             "@              	             �?���Q��?             @                          �]@�q�q�?             @������������������������       �                     �?                          �]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @       4                    �?\�sե��?A            �\@                           @D@d��4�o�?4            �W@������������������������       �                     $@       #                    �?�H�a��?/            @U@       "                    �J@`�Q��?             9@       !                   8q@���!pc�?             &@                            ]@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     ,@$       3       
             �?r�q��?$             N@%       (                   �_@��[�p�?            �G@&       '                   �[@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @)       ,                   `i@�?�'�@�?             C@*       +                   �b@���y4F�?
             3@������������������������       �                     .@������������������������       �                     @-       .                    �I@�}�+r��?             3@������������������������       �                     &@/       0                    o@      �?              @������������������������       �                     @1       2                    r@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     *@5       6                   �^@R���Q�?             4@������������������������       �                     $@7       8                    �J@�z�G��?             $@������������������������       �                     @������������������������       �                     @:       {                    �?�>4և��?�             l@;       Z                    @L@<����=�?z            �h@<       C                    �?�T�2�?\            �b@=       B                    �?�����H�?             ;@>       ?                   �g@H%u��?             9@������������������������       �        
             5@@       A                   �h@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @D       E                    �? @|���?O            �^@������������������������       �                     C@F       W                   `]@�8��8��?8             U@G       V                    �?���Q��?             .@H       O                    c@�	j*D�?             *@I       J                   �_@���Q��?             @������������������������       �                     �?K       L       	          �����      �?             @������������������������       �                     �?M       N                    @I@�q�q�?             @������������������������       �                      @������������������������       �                     �?P       U                   �p@      �?              @Q       T                    f@      �?             @R       S                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @X       Y                   `X@@	tbA@�?,            @Q@������������������������       �                     �?������������������������       �        +             Q@[       b                    �?~���L0�?            �H@\       a                   pb@      �?	             0@]       ^                    �?r�q��?             @������������������������       �                     @_       `                     @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@c       v                    �?4���C�?            �@@d       u       	          ����?��>4և�?             <@e       j                    �?� �	��?             9@f       g                   @`@X�<ݚ�?             "@������������������������       �                     @h       i       	          ����?�q�q�?             @������������������������       �                     @������������������������       �                      @k       t                    @      �?
             0@l       m                   �V@և���X�?	             ,@������������������������       �                      @n       o                   �m@�q�q�?             (@������������������������       �                     @p       q                     M@z�G�z�?             @������������������������       �                      @r       s                   ps@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @w       z                    a@���Q��?             @x       y                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?|       }                    `@�θ�?             :@������������������������       �                     @~       �                    b@���N8�?             5@       �       	          ����?      �?              @�       �                     L@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     *@�       �                    �?61���r�?�            Pv@�       �       	          ���@N1���?&            �N@�       �                    �?����3��?!             J@������������������������       �                     *@�       �                   �V@Hث3���?            �C@������������������������       �                     @�       �                   `c@j���� �?             A@�       �                   �Z@����X�?             <@�       �                   0r@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �E@�q�q�?             8@������������������������       �                     @�       �                   (q@�����?             5@������������������������       �                     .@�       �                    @O@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     "@�       �                    @E@P�0�e��?�            �r@�       �       	          033�?���Q��?             4@������������������������       �                     @�       �       
             �?�t����?             1@������������������������       �                     �?�       �                    �?      �?             0@�       �                    �?�8��8��?             (@������������������������       �                     $@�       �                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?�       �                   `_@�	��X�?�            @q@�       �                   �Q@���(-�?^            @b@�       �                   �l@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?@ݚ)�?\             b@�       �                    @H��2�?@            @W@�       �                    �?hl �&�??             W@�       �                   �s@�k~X��?.             R@������������������������       �        +            �P@�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �J@ףp=
�?             4@�       �                   q@r�q��?             @�       �                    @J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �]@@4և���?             ,@������������������������       �                     @�       �                    ^@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    \@���J��?            �I@�       �                   �[@`2U0*��?             9@������������������������       �        
             4@�       �                     R@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     :@�       �       	          ����?�N�#/�?S            @`@�       �       	          `ff�?�f7�z�?             =@�       �                    @K@r�q��?             @�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   0m@
;&����?             7@�       �                   �h@r�q��?             (@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                   �p@"pc�
�?             &@�       �                    �?�q�q�?             @������������������������       �                      @�       �                   @_@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                   �[@0�W���?B            @Y@�       �                    �?      �?             $@������������������������       �                      @�       �                   `@      �?              @������������������������       �                      @�       �                     K@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    n@H�g�}N�?;            �V@�       �                   @b@��s����?(            �O@�       �                   �m@PN��T'�?"             K@�       �                   �c@^�!~X�?!            �J@������������������������       �                    �B@�       �                    �N@     ��?             0@�       �                    _@      �?             (@�       �                   `l@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                    �?X�<ݚ�?             "@������������������������       �                      @�       �                   @d@����X�?             @�       �       	          `ff@���Q��?             @�       �                     L@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     <@q�tq�bh�h"h#K �q�h%�q�Rq�(KK�KK�q�hV�B�       �t@     y@     p@      ^@      P@     @V@      @     �A@      �?      <@      �?      $@              @      �?      @              �?      �?       @              �?      �?      �?      �?                      �?              2@       @      @       @      @       @      �?      �?              �?      �?      �?                      �?               @              @     �N@      K@      M@     �B@              $@      M@      ;@       @      1@       @      @       @      �?              �?       @                       @              ,@      I@      $@     �B@      $@      @      @      @                      @     �@@      @      .@      @      .@                      @      2@      �?      &@              @      �?      @              @      �?              �?      @              *@              @      1@              $@      @      @      @                      @      h@      ?@     �e@      9@     `a@      $@      8@      @      6@      @      5@              �?      @              @      �?               @             �\@      @      C@             @S@      @      "@      @      "@      @       @      @              �?       @       @      �?              �?       @               @      �?              @      �?      @      �?      �?      �?      �?                      �?       @              @                       @      Q@      �?              �?      Q@              A@      .@      .@      �?      @      �?      @               @      �?       @                      �?      $@              3@      ,@      1@      &@      ,@      &@      @      @              @      @       @      @                       @      $@      @       @      @               @       @      @      @              �?      @               @      �?       @      �?                       @       @              @               @      @      �?      @      �?                      @      �?              4@      @              @      4@      �?      @      �?      @      �?      @                      �?      @              *@              S@     �q@     �@@      <@     �@@      3@      *@              4@      3@              @      4@      ,@      4@       @      �?      @              @      �?              3@      @              @      3@       @      .@              @       @      @                       @              @              "@     �E@     �o@       @      (@      @              @      (@      �?              @      (@      �?      &@              $@      �?      �?      �?                      �?      @      �?      @                      �?     �A@      n@      @     �a@      �?      �?              �?      �?              @     `a@      @     @V@      @     @V@      �?     �Q@             �P@      �?      @              @      �?               @      2@      �?      @      �?      �?              �?      �?                      @      �?      *@              @      �?      @      �?                      @      �?              �?      I@      �?      8@              4@      �?      @              @      �?                      :@      =@     @Y@      (@      1@      �?      @      �?      �?              �?      �?                      @      &@      (@       @      $@       @       @               @       @                       @      "@       @      @       @       @               @       @       @                       @      @              1@      U@      @      @       @              @      @       @              �?      @      �?                      @      (@     �S@      (@     �I@       @      G@      @      G@             �B@      @      "@      @      "@      @      @      @                      @              @      @              �?              @      @       @               @      @       @      @       @       @               @       @                      �?               @              <@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJu�7hG        hNhG        h<Kh=Kh>h"h#K �q�h%�q�Rq�(KK�q�hV�C              �?q�tq�bhJhZhEC       q��q�Rq�h^Kh_h`Kh"h#K �q�h%�q�Rq�(KK�q�hE�C       q�tq�bK�q�Rq�}q�(hKhjMhkh"h#K �q�h%�q�Rq�(KM�q�hr�Bx=         �       	          ����?p�Vv���?�           ��@       #                    �?X~�pX��?�            �v@              
             �?���!���?3            �S@                           �L@      �?             (@������������������������       �                     @                          8r@���Q��?             @������������������������       �                      @������������������������       �                     @	                           �?�qM�R��?+            �P@
                           �?d}h���?	             ,@                           �D@8�Z$���?             *@������������������������       �                     �?              	          ����?�8��8��?             (@������������������������       �                      @              	            �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?                           �H@ �h�7W�?"            �J@������������������������       �                     @@                          @V@؇���X�?             5@                           @O@      �?              @������������������������       �                     �?������������������������       �                     �?                           [@�KM�]�?             3@                          @_@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �?      �?             0@������������������������       �                     $@                           �q@r�q��?             @������������������������       �                     @!       "                   @`@      �?              @������������������������       �                     �?������������������������       �                     �?$       a                    �?�9!���?�            �q@%       X                    �?4uj�w��?K            @\@&       S       
             �?,��I�?8            �U@'       8                    �H@P��E��?.             R@(       3                   �^@�������?             >@)       2                   �p@և���X�?	             ,@*       -       
             �?      �?              @+       ,                     G@      �?              @������������������������       �                     �?������������������������       �                     �?.       1                   pc@r�q��?             @/       0                   @b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @4       5                   �e@      �?	             0@������������������������       �                     *@6       7                    �D@�q�q�?             @������������������������       �                      @������������������������       �                     �?9       N                   �a@�G��l��?             E@:       E                   `_@���Q��?            �A@;       <                    �?X�Cc�?	             ,@������������������������       �                      @=       D                    �O@      �?             (@>       ?                   �`@"pc�
�?             &@������������������������       �                     @@       A                    W@�q�q�?             @������������������������       �                     @B       C                   0a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?F       G                   �b@���N8�?             5@������������������������       �                     (@H       I                   @`@X�<ݚ�?             "@������������������������       �                     @J       K                     L@z�G�z�?             @������������������������       �                      @L       M                   0a@�q�q�?             @������������������������       �                      @������������������������       �                     �?O       P                   �b@؇���X�?             @������������������������       �                     @Q       R                    �J@      �?             @������������������������       �                     �?������������������������       �                     @T       W                    �P@��S���?
             .@U       V                    T@�q�q�?	             (@������������������������       �                     @������������������������       �                      @������������������������       �                     @Y       Z       	          ����?8�Z$���?             :@������������������������       �                     0@[       `                     L@���Q��?             $@\       _       
             �?z�G�z�?             @]       ^                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @b       �                    @���PL6�?l            �e@c       l                   �X@�npº��?a            �b@d       e                   �j@���!pc�?	             &@������������������������       �                     @f       i                    �?և���X�?             @g       h                   �m@      �?              @������������������������       �                     �?������������������������       �                     �?j       k                    @I@���Q��?             @������������������������       �                      @������������������������       �                     @m       z                    �K@�d�g��?X            �a@n       w                   �g@������?C             [@o       v                   �a@�O4R���?A            �Z@p       q                    @B@ >�֕�?            �A@������������������������       �                     �?r       s                    �?г�wY;�?             A@������������������������       �                     @@t       u                   @^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        ,            �Q@x       y                    �D@      �?              @������������������������       �                     �?������������������������       �                     �?{       �                   �a@     ��?             @@|       �                    @M@�\��N��?             3@}       �                    �?�<ݚ�?             "@~                          @_@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �       	          ����?�z�G��?             $@�       �                    �?���Q��?             @������������������������       �                     �?�       �                   `Z@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     *@�       �                   �p@8�A�0��?             6@�       �                    �?���Q��?             .@�       �                   �d@���Q��?             $@�       �                   c@և���X�?             @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?�zц��?�            w@�       �                   �R@�'�=z��?&            �P@������������������������       �                     @�       �                     P@��S���?#             N@�       �                   �a@� �	��?             I@�       �       	          033�?X�<ݚ�?             B@�       �                    �C@���N8�?             5@������������������������       �                      @�       �                   �p@�S����?             3@������������������������       �                     (@�       �                   pb@և���X�?             @�       �                   @_@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    a@������?
             .@������������������������       �                     @�       �                   @n@X�<ݚ�?             "@������������������������       �                     @�       �                    �K@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �c@؇���X�?	             ,@�       �                   `c@$�q-�?             *@�       �       
             �?r�q��?             @������������������������       �                     @�       �                   pm@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�       �                   h@�DÓ ��?�            �r@�       �                    �?X'"7��?I             [@�       �                    @M@p�C��?<            �V@������������������������       �                     �H@�       �                   P`@���N8�?             E@�       �                    `@ ���J��?            �C@�       �                   `_@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     =@�       �                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @O@@�0�!��?             1@�       �                   �d@��S�ۿ?             .@������������������������       �        	             &@�       �                   �d@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�                         �b@8�f�ȭ�?�            `h@�       �                   �j@H�ՠ&��?o            @d@�       �                   �h@      �?             2@������������������������       �                      @�       �                   �j@     ��?             0@�       �                    �L@X�Cc�?             ,@�       �       
             �?����X�?             @�       �                    �G@���Q��?             @������������������������       �                      @�       �                    @L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�                          �P@�8��8��?b             b@�                           `P@����y7�?V            @_@�       �                   �v@85�}C�?T            �^@�       �       	          ����? ,��-�?R            �]@�       �       
             �?�d�����?             3@������������������������       �                     @�       �                    �N@�q�q�?             .@�       �                     M@      �?             $@�       �                    �?����X�?             @�       �                    �?r�q��?             @������������������������       �                     �?�       �                    �?z�G�z�?             @�       �                   �[@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �D@Pa�	�?C            �X@�       �       
             �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �? r���?@            �W@������������������������       �                     1@�       �                   �`@ ���J��?3            �S@�       �                    �N@�t����?             1@�       �                   po@$�q-�?             *@������������������������       �                     @�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?             @�       �       	          `ff�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �        %            �N@�       �                    �K@      �?             @������������������������       �                      @������������������������       �                      @            	          `ff�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     3@                        �[@�'�=z��?            �@@������������������������       �                      @                         @�g�y��?             ?@                         �?
j*D>�?             :@	            	             �?���|���?             &@
                        Pe@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @            	             @������?
             .@                         �?�8��8��?             (@                        Pd@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @                         �E@z�G�z�?             @                        �j@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @q�tq�bh�h"h#K �q�h%�q�Rq�(KMKK�q�hV�B�       @t@     �y@     @o@     �\@     �Q@      "@      "@      @      @               @      @       @                      @     �N@      @      &@      @      &@       @              �?      &@      �?       @              @      �?              �?      @                      �?      I@      @      @@              2@      @      �?      �?              �?      �?              1@       @       @      �?       @                      �?      .@      �?      $@              @      �?      @              �?      �?      �?                      �?     �f@     �Z@     �D@      R@     �B@      I@      =@     �E@      @      7@      @       @      @       @      �?      �?              �?      �?              @      �?      �?      �?      �?                      �?      @                      @      �?      .@              *@      �?       @               @      �?              6@      4@      5@      ,@      @      "@       @              @      "@       @      "@              @       @      @              @       @      �?       @                      �?      �?              0@      @      (@              @      @              @      @      �?       @               @      �?       @                      �?      �?      @              @      �?      @      �?                      @       @      @       @      @              @       @                      @      @      6@              0@      @      @      @      �?      �?      �?      �?                      �?      @                      @     `a@      A@     @`@      5@      @       @              @      @      @      �?      �?      �?                      �?       @      @       @                      @     �_@      *@     @Z@      @      Z@       @     �@@       @              �?     �@@      �?      @@              �?      �?              �?      �?             �Q@              �?      �?      �?                      �?      6@      $@      "@      $@       @      @       @       @               @       @                      @      @      @       @      @      �?              �?      @      �?                      @      @              *@              "@      *@      "@      @      @      @      @      @      �?      @              @      �?              @                      @      @                      @     �R@     pr@      @@      A@              @      @@      <@      6@      <@      4@      0@      0@      @               @      0@      @      (@              @      @      �?      @      �?                      @      @              @      &@              @      @      @      @              �?      @      �?                      @       @      (@      �?      (@      �?      @              @      �?      �?      �?                      �?              @      �?              $@              E@     Pp@      @     �Y@       @     @V@             �H@       @      D@      �?      C@      �?      "@              "@      �?                      =@      �?       @      �?                       @      @      ,@      �?      ,@              &@      �?      @              @      �?               @             �B@     �c@      5@     �a@      "@      "@       @              @      "@      @      "@      @       @      @       @       @              �?       @               @      �?               @                      @       @              (@     �`@      (@     @\@      $@      \@       @     �[@      @      ,@              @      @      $@      @      @       @      @      �?      @              �?      �?      @      �?      @      �?                      @              �?      �?              @                      @      @      X@      �?      @              @      �?               @     @W@              1@       @      S@       @      .@      �?      (@              @      �?      @              @      �?              �?      @      �?      �?      �?                      �?               @             �N@       @       @       @                       @       @      �?              �?       @                      3@      0@      1@               @      0@      .@      .@      &@      @      @      �?      @              @      �?              @              &@      @      &@      �?      @      �?              �?      @              @                      @      �?      @      �?      �?      �?                      �?              @q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ��!XhG        hNhG        h<Kh=Kh>h"h#K �q�h%�q�Rq�(KK�q�hV�C              �?q�tq�bhJhZhEC       qنq�Rq�h^Kh_h`Kh"h#K �q�h%�q�Rq�(KK�q�hE�C       q�tq�bK�q�Rq�}q�(hKhjMhkh"h#K �q�h%�q�Rq�(KM�q�hr�B=         �       	          ����?U�ք�?�           ��@       G                    �?��R�{�?�             w@                          @E@��\���?Z             a@                           [@�?�|�?            �B@       
                    �?@4և���?	             ,@       	                    �J@�����H�?             "@                           @G@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     7@       F                   �f@�eP*L��?D            �X@       ;       	          833�?I� ��?A             W@       6                    �?��J�fj�?4            �R@       5       
             �?      �?-             N@                          �`@j���� �?(            �I@                           �?؇���X�?             ,@������������������������       �                      @                           `@r�q��?	             (@������������������������       �                     @                            I@����X�?             @                          �l@      �?              @������������������������       �                     �?������������������������       �                     �?                          @h@z�G�z�?             @������������������������       �                     @������������������������       �                     �?       0                    �L@��+��?            �B@       '                    `@���Q��?             >@       &                    @K@     ��?             0@        !       
             �?X�Cc�?
             ,@������������������������       �                      @"       %                    ]@�q�q�?             (@#       $                   pd@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @(       )                    �D@d}h���?             ,@������������������������       �                     �?*       /                   c@8�Z$���?             *@+       ,                    �G@���Q��?             @������������������������       �                     �?-       .                   �m@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @1       4                   �l@؇���X�?             @2       3                   @d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     "@7       8                   �p@؇���X�?             ,@������������������������       �                     "@9       :                    @I@���Q��?             @������������������������       �                      @������������������������       �                     @<       E                   pd@r�q��?             2@=       D                    �?�t����?             1@>       C                    �L@      �?             0@?       B                   ``@r�q��?             @@       A                   `m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     $@������������������������       �                     �?������������������������       �                     �?������������������������       �                     @H       �                    @�'�f7��?�             m@I       N                    @H@�y�b�w�?�             k@J       K                    �?�|���?=             V@������������������������       �        :            �T@L       M                    V@r�q��?             @������������������������       �                     �?������������������������       �                     @O       �                   @g@     ��?T             `@P       S                   �Z@4�=ݍ�?S            �_@Q       R                   �`@      �?             @������������������������       �                     @������������������������       �                     @T       _                   @Z@��p��?O            @^@U       V                    @M@      �?
             (@������������������������       �                     @W       X                    �?�q�q�?             "@������������������������       �                     �?Y       ^                   �X@      �?              @Z       [                    �N@؇���X�?             @������������������������       �                     @\       ]                   �l@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?`       a                    �?����?E            @[@������������������������       �                    �E@b       �                   �e@j�'�=z�?'            �P@c       z       
             �?     ��?&             P@d       s       	          833�?�{��?��?             K@e       p                   @t@X�EQ]N�?            �E@f       i                   �`@��(\���?             D@g       h                   �_@�q�q�?             @������������������������       �                     @������������������������       �                      @j       k                   �q@г�wY;�?             A@������������������������       �                     =@l       o                    �?z�G�z�?             @m       n                    �L@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @q       r                   u@�q�q�?             @������������������������       �                      @������������������������       �                     �?t       u                   @i@�eP*L��?             &@������������������������       �                      @v       w                    _@�q�q�?             "@������������������������       �                      @x       y                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @{       �                   �m@���Q��?	             $@|       }                    �L@      �?              @������������������������       �                     @~                            P@z�G�z�?             @������������������������       �                     @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                   �c@     ��?
             0@�       �                   a@�eP*L��?             &@������������������������       �                     @�       �                   `Q@����X�?             @������������������������       �                     �?�       �                   �_@r�q��?             @�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�                           �?��@�yC�?�            �v@�       �                    @K@���mC�?�            �o@�       �                   q@��7Y��?I            �[@�       �       	             @rѱ�D��?:            �V@�       �                    �?��%��?.            �R@�       �                    �?�������?             A@�       �                    _@X�<ݚ�?             "@������������������������       �                     @�       �                    Z@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �m@�J�4�?             9@������������������������       �                     4@�       �                   `^@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �\@R���Q�?             D@������������������������       �                     @�       �                    �?�MI8d�?            �B@������������������������       �                     1@�       �                   �c@�z�G��?             4@�       �                    @      �?             (@�       �                    �?      �?              @������������������������       �                     �?�       �                    �F@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �B@@�0�!��?             1@������������������������       �                     �?�       �                   �Z@      �?             0@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       
             �?$�q-�?	             *@������������������������       �                     @�       �                    �?r�q��?             @�       �       	             @z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �`@R���Q�?             4@�       �                    �?�q�q�?             "@�       �                    c@      �?              @�       �                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             &@�       �                    �?�E���-�?\             b@�       �                    �Q@�7��d��?=             Y@�       �       
             �?�FVQ&�?<            �X@�       �                   �_@�}��L�?+            �R@�       �                    �L@      �?             @@�       �       	             �?$�q-�?             *@�       �       	          ����?؇���X�?             @������������������������       �                     @�       �                    @L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     3@������������������������       �                    �E@�       �                   �X@�q�q�?             8@������������������������       �                     �?�       �                    @M@�㙢�c�?             7@������������������������       �                     @�       �       	          ����?      �?             0@�       �                   �`@X�<ݚ�?             "@������������������������       �                     @�       �                    �M@r�q��?             @�       �       	             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    �O@���|���?             F@�       �                    �?<ݚ)�?             B@�       �                    �N@����X�?             @�       �                     @r�q��?             @�       �                   xu@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                   �r@V�a�� �?             =@�       �                   �e@�>4և��?             <@�       �                   �p@ȵHPS!�?             :@�       �       	          ����?���}<S�?             7@�       �                    �N@����X�?             @�       �                    @M@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     0@�       �                    �?�q�q�?             @������������������������       �                     �?�       �       	          `ff�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                     Q@      �?              @������������������������       �                     @�       �                   �a@      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                         �?���l��?E            �[@            	          033�?���7�?6             V@                        �x@ ��ʻ��?)             Q@������������������������       �        '            �P@                        ��@      �?              @������������������������       �                     �?������������������������       �                     �?      	                  `c@R���Q�?             4@������������������������       �                     "@
                        �r@���!pc�?             &@������������������������       �                      @������������������������       �                     @                         �?�㙢�c�?             7@                        pc@���!pc�?	             &@            	          ����?      �?              @������������������������       �                     �?������������������������       �                     @                         e@�q�q�?             @������������������������       �                      @������������������������       �                     �?                        p`@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@q�tq�bh�h"h#K �q�h%�q�Rq�(KMKK�q�hV�Bp        t@     �y@     �n@     �^@     �K@     @T@      �?      B@      �?      *@      �?       @      �?      �?              �?      �?                      @              @              7@      K@     �F@     �G@     �F@      @@      E@      >@      >@      5@      >@       @      (@               @       @      $@              @       @      @      �?      �?              �?      �?              �?      @              @      �?              3@      2@      2@      (@      @      "@      @      "@               @      @      @      @       @      @                       @              @       @              &@      @              �?      &@       @      @       @              �?      @      �?      @                      �?       @              �?      @      �?      �?              �?      �?                      @      "@               @      (@              "@       @      @       @                      @      .@      @      .@       @      .@      �?      @      �?      �?      �?      �?                      �?      @              $@                      �?              �?      @             �g@      E@      g@      ?@     �U@      �?     �T@              @      �?              �?      @             �X@      >@     �X@      =@      @      @              @      @             �W@      :@      @      "@              @      @      @      �?               @      @      �?      @              @      �?      @      �?                      @      �?              W@      1@     �E@             �H@      1@     �H@      .@     �E@      &@      C@      @     �B@      @      @       @      @                       @     �@@      �?      =@              @      �?       @      �?              �?       @               @              �?       @               @      �?              @      @       @              @      @       @              �?      @      �?                      @      @      @      @      @      @              �?      @              @      �?      �?      �?                      �?       @                       @              �?      @      &@      @      @              @      @       @              �?      @      �?       @      �?       @                      �?      @                      @     @S@     r@     @Q@     @g@      G@     @P@     �E@      H@      D@      A@      "@      9@      @      @              @      @      �?              �?      @              @      5@              4@      @      �?              �?      @              ?@      "@              @      ?@      @      1@              ,@      @      @      @       @      @              �?       @      @       @                      @      @               @              @      ,@      �?               @      ,@      �?       @      �?                       @      �?      (@              @      �?      @      �?      @      �?                      @              �?      @      1@      @      @       @      @      �?      @      �?                      @      �?              �?                      &@      7@     @^@      @     @W@      @     @W@      �?     �R@      �?      ?@      �?      (@      �?      @              @      �?      �?              �?      �?                      @              3@             �E@      @      3@      �?              @      3@              @      @      (@      @      @      @              �?      @      �?      @              @      �?                       @              @      �?              0@      <@      &@      9@      @       @      @      �?      @      �?      @                      �?       @                      �?      @      7@      @      7@      @      7@       @      5@       @      @       @       @               @       @                      @              0@      �?       @              �?      �?      �?      �?                      �?       @              �?              @      @      @              �?      @      �?      �?              �?      �?                       @       @     �Y@      @      U@      �?     �P@             �P@      �?      �?      �?                      �?      @      1@              "@      @       @               @      @              @      3@      @       @      �?      @      �?                      @       @      �?       @                      �?      �?      &@      �?                      &@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJC�NhG        hNhG        h<Kh=Kh>h"h#K �q�h%�q�Rq�(KK�q�hV�C              �?q�tq�bhJhZhEC       q��q�Rq�h^Kh_h`Kh"h#K �q�h%�q�Rq�(KK�q�hE�C       r   tr  bK�r  Rr  }r  (hKhjMhkh"h#K �r  h%�r  Rr  (KM�r  hr�B�>         �                    �?4�5����?�           ��@       �                    �?����&�?           Py@       2                   `_@Ј�^�i�?�            @r@                           �?֦:O���?X             b@              	          ����?��<D�m�??            �X@                           �O@�r����?             >@              	          hff�?ܷ��?��?             =@                          @W@`2U0*��?             9@	       
                    @I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     7@                          �\@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?                           _@г�wY;�?-             Q@                           �?0�z��?�?(             O@              
             �?r�q��?             @������������������������       �                      @                           �H@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        %             L@                          �[@r�q��?             @������������������������       �                     @              	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?       -                   �q@֭��F?�?            �G@       $       	          @33�?      �?             A@        #                   �Z@@4և���?             ,@!       "       	             �z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@%       ,                     M@z�G�z�?	             4@&       '                   �W@�q�q�?             (@������������������������       �                     @(       )                   Pk@�q�q�?             @������������������������       �                     @*       +                    a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @.       1                   �r@$�q-�?             *@/       0       	             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@3       p       	          ����?|���?e            `b@4       g                   Pd@�xGZ���?G            @Z@5       D       
             �?X��ʑ��?:            �U@6       ?       	            �?�z�G��?             4@7       :                   c@X�Cc�?
             ,@8       9                   �a@      �?             @������������������������       �                     @������������������������       �                     �?;       >                    �?z�G�z�?             $@<       =                    @M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @@       A                    c@r�q��?             @������������������������       �                     @B       C                   @_@�q�q�?             @������������������������       �                      @������������������������       �                     �?E       F                    @C@�eP*L��?+            �P@������������������������       �                     @G       \                   Pb@Ɣ��Hr�?&            �M@H       K                    �?�X���?             F@I       J                    a@      �?             $@������������������������       �                     @������������������������       �                     @L       M                   �^@�t����?             A@������������������������       �                     (@N       S                   �j@�eP*L��?             6@O       P       	          ����?�z�G��?             $@������������������������       �                     @Q       R       	             �?      �?             @������������������������       �                     @������������������������       �                     �?T       Y                   �`@�q�q�?             (@U       X                    `@      �?              @V       W                   �b@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @Z       [                   Xp@      �?             @������������������������       �                     �?������������������������       �                     @]       f                    �?��S���?             .@^       a                    �J@�n_Y�K�?
             *@_       `                    d@      �?              @������������������������       �                     @������������������������       �                     �?b       c                   d@z�G�z�?             @������������������������       �                     @d       e                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @h       k                    �?���y4F�?             3@i       j                   pf@      �?              @������������������������       �                     @������������������������       �                     @l       o                    �D@�C��2(�?             &@m       n                    a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@q       r                   �`@�����?             E@������������������������       �                     "@s       t                   @M@<���D�?            �@@������������������������       �                     �?u       ~                    �?     ��?             @@v       w                    �?"pc�
�?             &@������������������������       �                     @x       y                     J@���Q��?             @������������������������       �                     �?z       {                   0k@      �?             @������������������������       �                      @|       }                   `a@      �?              @������������������������       �                     �?������������������������       �                     �?       �                   @a@���N8�?             5@������������������������       �                     &@�       �                   �p@ףp=
�?             $@������������������������       �                      @�       �                   pd@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       
             �?h��)�~�?K            @\@�       �                   �Q@<���D�?1            �P@������������������������       �                      @�       �                    `R@     ��?0             P@�       �                    �?�[|x��?/            �O@�       �                    �?�����H�?             "@�       �                   0n@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �a@�>����?)             K@�       �                    _@ qP��B�?"            �E@������������������������       �                     ;@�       �       	             �?      �?             0@�       �                   �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     *@�       �                     K@���!pc�?             &@�       �       	          833�?և���X�?             @�       �                   �c@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                   �`@=QcG��?            �G@������������������������       �                    �@@�       �                     J@d}h���?             ,@�       �                   �b@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�       �                    �K@������?�            �t@�       �                   �g@��UTF@�?�            @k@�       �       	          ����?�ӭ�a��?�             k@�       �                    �?�7��?f            �c@�       �                    �J@ pƵHP�?             J@������������������������       �                    �F@�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �       
             �?�q-�?G             Z@�       �                   �a@$�q-�?>            �V@�       �                    �?PN��T'�?             ;@������������������������       �                     �?�       �                    �B@8�Z$���?             :@������������������������       �                     @�       �                   �Z@�nkK�?             7@�       �                    @I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     5@�       �                   @[@     �?,             P@�       �                    �H@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   `]@�g�y��?*             O@�       �                   p@      �?              @������������������������       �                     @�       �                    \@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       
             �?@3����?%             K@������������������������       �                     $@�       �                    @`���i��?             F@������������������������       �                    �E@������������������������       �                     �?������������������������       �        	             *@�       �       
             �?�q�q�?&             N@������������������������       �                     &@�       �                    �?�`���?!            �H@�       �       	             @�eP*L��?             F@�       �                    �?^H���+�?            �B@�       �                    �?8�Z$���?
             *@������������������������       �                     @�       �                   `d@����X�?             @������������������������       �                     @�       �                   0e@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   @^@r�q��?             8@�       �       	          ����?�C��2(�?             &@�       �                    ]@؇���X�?             @������������������������       �                     @�       �                   �b@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �c@�θ�?             *@������������������������       �                     @�       �                    @      �?             @�       �                    q@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �?��+��?N            �[@�       �       	          ����?��X��?             <@�       �                    _@؇���X�?             5@�       �                   �Z@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �c@      �?             0@������������������������       �                     ,@�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �L@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?F~��7�?6            �T@�       �                    �Q@�����?             5@�       �       	          ����?P���Q�?             4@������������������������       �                     ,@�       �                   `Z@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�             	          ����?r֛w���?(             O@             	          ����?     ��?             @@                          Q@�	j*D�?             :@                        �d@      �?             8@                        �d@��<b���?             7@                         �?�KM�]�?             3@                        pk@z�G�z�?             $@������������������������       �                     @      
      
             �?�q�q�?             @      	                   _@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@                        �c@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                         _@r�q��?             @                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                         @O@ףp=
�?             >@������������������������       �        
             0@                          P@d}h���?             ,@������������������������       �                     �?                         @R@8�Z$���?             *@                        �[@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @r	  tr
  bh�h"h#K �r  h%�r  Rr  (KMKK�r  hV�B�       �t@     y@      X@     Ps@     @U@     �i@      8@     @^@      @      W@      @      :@      @      :@      �?      8@      �?      �?      �?                      �?              7@       @       @       @                       @      �?               @     �P@      �?     �N@      �?      @               @      �?      @              @      �?                      L@      �?      @              @      �?      �?              �?      �?              2@      =@      1@      1@      *@      �?      @      �?              �?      @              "@              @      0@      @       @              @      @       @      @              �?       @      �?                       @               @      �?      (@      �?      @      �?                      @              "@     �N@     �U@     �L@      H@      E@      F@      @      ,@      @      "@      @      �?      @                      �?       @       @       @      �?       @                      �?              @      �?      @              @      �?       @               @      �?              B@      >@              @      B@      7@      =@      .@      @      @      @                      @      8@      $@      (@              (@      $@      @      @      @              �?      @              @      �?              @      @       @      @       @       @       @                       @              @      @      �?              �?      @              @       @      @       @      �?      @              @      �?              @      �?      @              �?      �?      �?                      �?       @              .@      @      @      @              @      @              $@      �?      �?      �?      �?                      �?      "@              @      C@              "@      @      =@      �?              @      =@       @      "@              @       @      @      �?              �?      @               @      �?      �?      �?                      �?      �?      4@              &@      �?      "@               @      �?      �?      �?                      �?      &@     �Y@       @      M@       @              @      M@      @      M@      �?       @      �?      �?              �?      �?                      @      @      I@      �?      E@              ;@      �?      .@      �?       @               @      �?                      *@      @       @      @      @      @      �?      @                      �?              @              @      �?              @      F@             �@@      @      &@      @      �?      @                      �?              $@     �m@      W@     �f@     �A@     �f@     �@@     �b@       @     �I@      �?     �F@              @      �?      @                      �?     @X@      @      U@      @      7@      @      �?              6@      @              @      6@      �?      �?      �?      �?                      �?      5@             �N@      @      �?      �?              �?      �?              N@       @      @      �?      @              �?      �?      �?                      �?     �J@      �?      $@             �E@      �?     �E@                      �?      *@             �A@      9@      &@              8@      9@      8@      4@      8@      *@      &@       @      @              @       @      @              �?       @               @      �?              *@      &@      $@      �?      @      �?      @              @      �?              �?      @              @              @      $@              @      @      @       @      @              @       @              �?                      @              @               @      K@     �L@      3@      "@      2@      @      @       @               @      @              .@      �?      ,@              �?      �?              �?      �?              �?      @      �?                      @     �A@      H@      3@       @      3@      �?      ,@              @      �?              �?      @                      �?      0@      G@      *@      3@       @      2@      @      2@      @      2@       @      1@       @       @              @       @      @       @      �?       @                      �?              @              "@      @      �?      @                      �?      �?               @              @      �?      �?      �?              �?      �?              @              @      ;@              0@      @      &@      �?               @      &@       @      @       @                      @              @r  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJ�R�[hG        hNhG        h<Kh=Kh>h"h#K �r  h%�r  Rr  (KK�r  hV�C              �?r  tr  bhJhZhEC       r  �r  Rr  h^Kh_h`Kh"h#K �r  h%�r  Rr  (KK�r  hE�C       r   tr!  bK�r"  Rr#  }r$  (hKhjK�hkh"h#K �r%  h%�r&  Rr'  (KK��r(  hr�Bx6         �       	          ����?6������?�           ��@       u                    �?��_���?�             w@       6                    �?�������?�             s@       -                    �?�G��l��?B            @Z@       "                   xp@��6���?7             U@                            E@��۾%d�?)             M@                           �?؇���X�?             @������������������������       �                     �?	       
                   �\@r�q��?             @������������������������       �                     @                           a@�q�q�?             @������������������������       �                     �?������������������������       �                      @       !                   `c@�"U����?$            �I@                          @E@�q�q�?"             H@������������������������       �                     @                          �_@�%^�?            �E@                          �l@���|���?	             &@              
             �?      �?              @                           �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                          pi@      �?             @@                          �b@�θ�?
             *@������������������������       �                     $@������������������������       �                     @               
             �?�}�+r��?             3@                           �L@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     ,@������������������������       �                     @#       &                    �?���B���?             :@$       %                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @'       (                    `@���N8�?
             5@������������������������       �                     (@)       *                   8r@�����H�?             "@������������������������       �                     @+       ,                   �`@      �?             @������������������������       �                     �?������������������������       �                     @.       3                   �`@��s����?             5@/       0       	            �?�����H�?	             2@������������������������       �                     (@1       2                    �M@�q�q�?             @������������������������       �                      @������������������������       �                     @4       5                     P@�q�q�?             @������������������������       �                     �?������������������������       �                      @7       T                    @L@�i'tU��?�             i@8       9                   `X@��e3���?e            �c@������������������������       �                     @:       I                   `]@��F��?d            `c@;       H                   �p@R�}e�.�?             :@<       =                    �?��Q��?             4@������������������������       �                     @>       ?                     G@      �?             ,@������������������������       �                     @@       G                    �J@���|���?             &@A       F                   �d@�<ݚ�?             "@B       C                   �X@���Q��?             @������������������������       �                     �?D       E                   @[@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @J       K                    �?�7�	|��?T             `@������������������������       �                    �C@L       M                    @K@�E�����?8            �V@������������������������       �        0            �S@N       S                    �K@�8��8��?             (@O       R       	          ����?z�G�z�?             @P       Q                   �n@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @U       `                    �?v ��?            �E@V       [       
             �?�t����?             1@W       X                   0o@      �?             @������������������������       �                     �?Y       Z       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?\       _                     P@�θ�?             *@]       ^                   �_@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@������������������������       �                      @a       j                    _@
j*D>�?             :@b       c                   �T@      �?              @������������������������       �                     �?d       e                    W@؇���X�?             @������������������������       �                     @f       i                    �?      �?             @g       h                    `@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?k       l                    �?�E��ӭ�?             2@������������������������       �                     @m       r                    @O@�n_Y�K�?	             *@n       q                    @�q�q�?             @o       p                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @s       t       	          ����?؇���X�?             @������������������������       �                     @������������������������       �                     �?v       w                    V@���@M^�?&             O@������������������������       �                     8@x       �       	          ����?p�ݯ��?             C@y       z       
             �?">�֕�?            �A@������������������������       �                      @{       �                     P@�5��?             ;@|       }                    [@�<ݚ�?             2@������������������������       �                      @~                           �?      �?             0@������������������������       �                     �?�       �                   �c@��S�ۿ?
             .@������������������������       �                     $@�       �                    @I@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    �Q@�<ݚ�?             "@�       �                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?xƅd�?�            �v@�       �                    f@`U���H�?�            �n@�       �                   �U@�R����?�            @n@������������������������       �                     �?�       �                   {@X{����?�             n@�       �                   �_@H�4�l��?�            �m@�       �                   `_@r�q��?-            �S@�       �                    �?$�Z����?,             S@�       �                   �j@�����H�?&            �O@�       �                   �i@"pc�
�?            �@@�       �                   �^@��� ��?             ?@������������������������       �                     (@�       �                     K@���y4F�?             3@������������������������       �                     *@�       �                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                   �s@(;L]n�?             >@������������������������       �                     ;@�       �                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @[@�	j*D�?             *@������������������������       �                     @�       �       	             @      �?              @�       �                   �n@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   @l@x�@�E-�?j             d@�       �                    �?�|���?6             V@������������������������       �        "            �J@�       �                    �?��?^�k�?            �A@�       �       	          ����?�IєX�?             1@�       �       	          033�?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@������������������������       �        	             2@�       �                   �l@����1�?4            @R@�       �                   �a@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   q@�IєX�?0             Q@������������������������       �                     =@�       �       	          ����?��-�=��?            �C@�       �                    �?      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �a@ >�֕�?            �A@�       �       	          033�?�KM�]�?             3@������������������������       �        
             *@�       �                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     0@������������������������       �                      @�       �                   �f@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �`@z���p��?G            @^@�       �                    �?��r._�?            �D@�       �       	          pff�?���Q��?             @������������������������       �                      @�       �                   `Z@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       
             �?�����H�?             B@�       �                   �n@      �?              @�       �                   @]@և���X�?             @������������������������       �                      @�       �                    �J@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �?h�����?             <@�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     :@�       �                    ]@��Q���?0             T@�       �                    f@�q�q�?             (@�       �                    @�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   Pe@��M���?*             Q@�       �       	          `ff@^l��[B�?#             M@�       �       	          ����?�t����?            �I@�       �                    d@���Q��?             @������������������������       �                     @������������������������       �                      @�       �       	          033�?���}<S�?             G@������������������������       �                     =@�       �                   �n@������?             1@������������������������       �        	             &@�       �                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �E@���Q��?             $@������������������������       �                      @�       �                    �?      �?              @������������������������       �                      @������������������������       �                     @r)  tr*  bh�h"h#K �r+  h%�r,  Rr-  (KK�KK�r.  hV�B�       �t@     �x@      o@     �]@      l@     @T@     �K@      I@      C@      G@     �@@      9@      �?      @              �?      �?      @              @      �?       @      �?                       @      @@      3@      @@      0@              @      @@      &@      @      @      �?      @      �?       @               @      �?                      @      @              <@      @      $@      @      $@                      @      2@      �?      @      �?      @                      �?      ,@                      @      @      5@      @      �?              �?      @              �?      4@              (@      �?       @              @      �?      @      �?                      @      1@      @      0@       @      (@              @       @               @      @              �?       @      �?                       @     @e@      ?@     `b@      &@              @     `b@       @      3@      @      *@      @      @              @      @      @              @      @       @      @       @      @      �?              �?      @              @      �?                      @       @              @              `@      �?     �C@             @V@      �?     �S@              &@      �?      @      �?      �?      �?      �?                      �?      @              @              7@      4@      (@      @       @       @      �?              �?       @               @      �?              $@      @      $@      �?              �?      $@                       @      &@      .@      @       @              �?      @      �?      @              @      �?       @      �?              �?       @              �?              @      *@              @      @       @      @       @      �?       @               @      �?              @              �?      @              @      �?              8@      C@              8@      8@      ,@      8@      &@       @              0@      &@      ,@      @               @      ,@       @              �?      ,@      �?      $@              @      �?              �?      @               @      @       @      @       @                      @              @              @     �U@     �q@      :@     `k@      8@     @k@      �?              7@     @k@      5@     @k@      *@     @P@      &@     @P@      @      L@      @      ;@      @      ;@              (@      @      .@              *@      @       @      @                       @       @              �?      =@              ;@      �?       @      �?                       @      @      "@              @      @      @      �?      @      �?                      @      @               @               @      c@      �?     �U@             �J@      �?      A@      �?      0@      �?      @              @      �?                      $@              2@      @     �P@      @       @      @                       @      @      P@              =@      @     �A@       @       @      �?      �?              �?      �?              �?      �?              �?      �?               @     �@@       @      1@              *@       @      @       @                      @              0@       @               @      �?       @                      �?      N@     �N@      @      A@      @       @       @              �?       @               @      �?              @      @@      @      @      @      @       @              �?      @      �?                      @              �?      �?      ;@      �?      �?      �?                      �?              :@     �J@      ;@      @       @      �?       @               @      �?              @             �H@      3@     �F@      *@     �F@      @      @       @      @                       @      E@      @      =@              *@      @      &@               @      @              @       @                      @      @      @       @               @      @       @                      @r/  tr0  bubhhubh)�r1  }r2  (hhh	h
hNhKhKhG        hh hNhJ�v}hG        hNhG        h<Kh=Kh>h"h#K �r3  h%�r4  Rr5  (KK�r6  hV�C              �?r7  tr8  bhJhZhEC       r9  �r:  Rr;  h^Kh_h`Kh"h#K �r<  h%�r=  Rr>  (KK�r?  hE�C       r@  trA  bK�rB  RrC  }rD  (hKhjM	hkh"h#K �rE  h%�rF  RrG  (KM	�rH  hr�B�9         �                    �?U�ք�?�           ��@       C       	          ����?r=ά�{�?�            Px@       
                    P@p�N�r�?_            �b@       	                    �D@      �?             @@                           �?      �?              @                          �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     8@                           _@4ʟ����?H            �]@                           �?�㙢�c�?             7@                           �?������?
             .@                           �O@8�Z$���?             *@                           �J@�8��8��?             (@������������������������       �                     @                           �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @       "                    �?�q�q��?:             X@                          �b@�㙢�c�?             7@                           �?�X�<ݺ?             2@������������������������       �        
             0@                          �o@      �?              @������������������������       �                     �?������������������������       �                     �?       !                   �c@���Q��?             @                            �N@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @#       0                   �b@�6����?+            @R@$       +                    �M@V������?            �B@%       &                    �?H%u��?             9@������������������������       �                     �?'       *                    �?�8��8��?             8@(       )                   �x@�r����?             .@������������������������       �        	             *@������������������������       �                      @������������������������       �                     "@,       /                    �?�q�q�?             (@-       .                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @1       B                    �?*O���?             B@2       A                   hp@�!���?             A@3       6                    �D@�G��l��?             5@4       5                    �B@z�G�z�?             @������������������������       �                     �?������������������������       �                     @7       8                    �E@      �?             0@������������������������       �                      @9       :                    \@և���X�?	             ,@������������������������       �                     @;       <                    �?z�G�z�?             $@������������������������       �                     @=       >                   0a@���Q��?             @������������������������       �                      @?       @                   �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �                      @D       E                   �U@��|Io��?�            �m@������������������������       �                     @F       Y                    �?0��x�-�?�            `m@G       H                    Y@д>��C�?             =@������������������������       �                      @I       X                    �?�����H�?             ;@J       W                   @e@R���Q�?             4@K       V                    �J@�KM�]�?             3@L       U       	             �?      �?              @M       T                    �?�q�q�?             @N       O                   @[@���Q��?             @������������������������       �                      @P       S       	             �?�q�q�?             @Q       R                    @I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     &@������������������������       �                     �?������������������������       �                     @Z       {                    �?p�eU}�?�            �i@[       j                   P`@T�n��?W             b@\       i                   �i@p� V�?;            �Y@]       ^                    @L@���7�?             F@������������������������       �        	             3@_       b                    �L@HP�s��?             9@`       a       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?c       d                    �?�nkK�?             7@������������������������       �                     &@e       h                    S@�8��8��?             (@f       g                   p`@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        %            �M@k       n                   @M@��P���?            �D@l       m                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @o       v       	          ����?(N:!���?            �A@p       q                   �a@      �?             @������������������������       �                     �?r       s                    \@���Q��?             @������������������������       �                      @t       u       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @w       z                   `j@XB���?             =@x       y       	          033@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     2@|       �                    �?0�z��?�?)             O@}       ~                   �r@`���i��?             F@������������������������       �                     D@       �                   `t@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     2@�       �                    I@ �>�?�            �u@�       �                   �]@���@��?            �B@�       �       
             �?�IєX�?
             1@�       �                   �\@      �?              @������������������������       �                     @�       �                   Pb@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                   `^@��Q��?             4@�       �                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �?d}h���?
             ,@������������������������       �                     �?�       �                    �G@�θ�?	             *@������������������������       �                     �?�       �                    �M@r�q��?             (@������������������������       �                     @�       �       	          `ff�?����X�?             @������������������������       �                     @�       �                   �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       	          ����?      �?�            @s@�       �                   �d@д>��C�?�             m@�       �                    [@t�6Z���?�            �k@�       �                    @N@���!pc�?             &@�       �                   �m@���Q��?             @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    @I@��^Oy�?�             j@�       �                    �?bۘ�W^�?L            @Z@�       �                   �c@��hJ,�?J            �Y@�       �                   �b@և���X�?             @������������������������       �                     @������������������������       �                     @�       �       	          ����?�W�{�5�?G            �W@�       �                    @���(`�?A            �U@�       �                    @G@@4և���??             U@�       �                   �a@0�z��?�?.             O@�       �                    �B@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        )            �K@�       �                   n@�GN�z�?             6@������������������������       �                     "@�       �                   `]@�n_Y�K�?	             *@������������������������       �                     @�       �                    �?�����H�?             "@�       �                   �q@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �[@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       
             �?      �?              @������������������������       �                      @�       �                   �j@      �?             @������������������������       �                      @�       �       	          ����?      �?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                   0a@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �^@�q-�?>             Z@������������������������       �                     ;@�       �                    �?�C��2(�?0            @S@������������������������       �                     ?@�       �                   Pj@*
;&���?             G@������������������������       �                     2@�       �       
             �?      �?             <@�       �                   �b@���B���?             :@�       �                    �K@      �?             4@������������������������       �                     �?�       �       
             �?���y4F�?             3@�       �                   a@      �?             @������������������������       �                      @������������������������       �                      @�       �                    _@�r����?	             .@������������������������       �                     �?�       �                    `P@@4և���?             ,@������������������������       �                     *@������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �       	          ����?�q�q�?             (@�       �                   �g@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   �`@:W��S��?*             S@�       �       
             �?�X���?             F@�       �                   �`@�n_Y�K�?            �C@�       �                    @P@      �?              @������������������������       �                     @������������������������       �                     �?�       �                    @B@r֛w���?             ?@������������������������       �                     �?�       �                   @_@�������?             >@�       �                    @�q�q�?             .@�       �                    j@      �?             $@������������������������       �                      @�       �                     H@      �?              @������������������������       �                     @�       �       
             �?���Q��?             @�       �       	          033�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �       	          `ff@�r����?             .@������������������������       �                     (@�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�                          �?     ��?             @@             
             �?�q�q�?             .@                        `c@r�q��?             (@                         �?�C��2(�?             &@������������������������       �                      @                        Pl@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     1@rI  trJ  bh�h"h#K �rK  h%�rL  RrM  (KM	KK�rN  hV�B�        t@     �y@     �T@      s@     �O@      V@      �?      ?@      �?      @      �?       @      �?                       @              @              8@      O@     �L@      @      3@      @      &@       @      &@      �?      &@              @      �?      @      �?                      @      �?               @                       @      M@      C@      3@      @      1@      �?      0@              �?      �?      �?                      �?       @      @       @      �?              �?       @                       @     �C@      A@      :@      &@      6@      @              �?      6@       @      *@       @      *@                       @      "@              @       @      @      �?              �?      @                      @      *@      7@      &@      7@      &@      $@      �?      @      �?                      @      $@      @       @               @      @              @       @       @      @              @       @       @              �?       @      �?                       @              *@       @              4@     @k@      @              1@     @k@      @      8@       @              @      8@      @      1@       @      1@       @      @       @      @       @      @               @       @      �?      �?      �?      �?                      �?      �?                      �?               @              &@      �?                      @      (@     @h@      &@     �`@       @     @Y@       @      E@              3@       @      7@      �?      �?              �?      �?              �?      6@              &@      �?      &@      �?      @      �?                      @              @             �M@      "@      @@      @      �?              �?      @              @      ?@      @      @      �?               @      @               @       @      �?              �?       @              �?      <@      �?      $@              $@      �?                      2@      �?     �N@      �?     �E@              D@      �?      @      �?                      @              2@     �m@     �Z@       @      =@      �?      0@      �?      @              @      �?      �?      �?                      �?              "@      @      *@      @       @      @                       @      @      &@              �?      @      $@      �?               @      $@              @       @      @              @       @      �?              �?       @             �l@     @S@      h@      D@     �g@      @@      @       @      @       @       @              �?       @      �?                       @              @      g@      8@      V@      1@     �U@      .@      @      @      @                      @      U@      &@     �S@       @     �S@      @     �N@      �?      @      �?              �?      @             �K@              1@      @      "@               @      @              @       @      �?      @      �?      @                      �?      @              �?       @      �?                       @      @      @       @              @      @       @              �?      @      �?       @      �?                       @              �?      �?       @               @      �?             @X@      @      ;@             �Q@      @      ?@             �C@      @      2@              5@      @      5@      @      .@      @              �?      .@      @       @       @       @                       @      *@       @              �?      *@      �?      *@                      �?      @                       @      @       @      @      @      @                      @              @     �C@     �B@      =@      .@      8@      .@      �?      @              @      �?              7@       @              �?      7@      @      $@      @      @      @               @      @      @      @               @      @       @      �?       @                      �?               @      @              *@       @      (@              �?       @      �?                       @      @              $@      6@      $@      @      $@       @      $@      �?       @               @      �?       @                      �?              �?              @              1@rO  trP  bubhhubh)�rQ  }rR  (hhh	h
hNhKhKhG        hh hNhJg}�XhG        hNhG        h<Kh=Kh>h"h#K �rS  h%�rT  RrU  (KK�rV  hV�C              �?rW  trX  bhJhZhEC       rY  �rZ  Rr[  h^Kh_h`Kh"h#K �r\  h%�r]  Rr^  (KK�r_  hE�C       r`  tra  bK�rb  Rrc  }rd  (hKhjK�hkh"h#K �re  h%�rf  Rrg  (KK��rh  hr�B�6         �                   �a@0����?�           ��@       )                   p`@�#V���?g           ��@       $                    �?�e/
�?G             [@                           �?������?&            �I@              	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @              	            �?�q�q�?$             H@	       
                   �\@���|���?             6@������������������������       �                      @              	          ����?�z�G��?             4@                          �^@@�0�!��?
             1@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                           I@�r����?             .@                           �?@4և���?             ,@                           `@ףp=
�?             $@                          �_@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @       !       
             �?$�q-�?             :@                          P`@�}�+r��?             3@������������������������       �                     .@                           @_@      �?             @              	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @"       #                    �N@؇���X�?             @������������������������       �                     @������������������������       �                     �?%       &                   �c@0�)AU��?!            �L@������������������������       �                     F@'       (       	          `ff@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?*       q                    �?~]@=���?            P|@+       L       	          ����?���Y)�?}            �i@,       ;                   �_@�K��&�?3            �U@-       :                    q@��
ц��?             J@.       9                    �?p�ݯ��?             C@/       4                   �i@">�֕�?            �A@0       1                    �?�����H�?             "@������������������������       �                     �?2       3       	          ����?      �?              @������������������������       �                     @������������������������       �                     �?5       8                    `@ȵHPS!�?             :@6       7                   �\@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �        	             2@������������������������       �                     @������������������������       �                     ,@<       I                    �?������?             A@=       H       	            �?r�q��?             >@>       ?       
             �?��<b���?             7@������������������������       �                     @@       A                    `@     ��?
             0@������������������������       �                     �?B       C                   �d@������?	             .@������������������������       �                     @D       G       
             �?�8��8��?             (@E       F                    �?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@������������������������       �                     �?������������������������       �                     @J       K                   �`@      �?             @������������������������       �                     @������������������������       �                     �?M       N                   �Q@؇���X�?J            �]@������������������������       �                      @O       Z                    �?�ݜ�?I            @]@P       Q                   h@���Q��?
             .@������������������������       �                     @R       W                     N@      �?             (@S       V                    ^@�����H�?             "@T       U       	             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @X       Y                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @[       j                    �?l��\��??            �Y@\       _                    �F@xdQ�m��?2            @T@]       ^                    @F@�r����?	             .@������������������������       �                     *@������������������������       �                      @`       c                   @i@���7�?)            �P@a       b       	          033�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?d       e                   �b@�]0��<�?&            �N@������������������������       �                     �I@f       g                    �?z�G�z�?             $@������������������������       �                     @h       i                    �J@����X�?             @������������������������       �                     @������������������������       �                      @k       p                    @M@��s����?             5@l       m                   �[@X�<ݚ�?             "@������������������������       �                      @n       o                    @J@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     (@r       �                    �?�A�9(��?�             o@s       t                    �?`-�I�w�?3             S@������������������������       �                     >@u       �       
             �?�q��/��?             G@v       y                   `X@�:�^���?            �F@w       x                   @_@�q�q�?             @������������������������       �                      @������������������������       �                     �?z       �                    �?@4և���?             E@{       |       
             �?P�Lt�<�?             C@������������������������       �                     *@}       ~                   �`@`2U0*��?             9@������������������������       �                     7@       �                   0b@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   @q@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �       	          ����?�������?p            �e@�       �                    ]@����l��?W             a@�       �       
             �?b�2�tk�?             2@������������������������       �                     �?�       �                   0f@j���� �?             1@�       �       	          ����?�q�q�?	             (@�       �                   `l@X�<ݚ�?             "@������������������������       �                     @�       �                   �p@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    @�D�d@6�?J            �]@�       �       	            �?,Z0R�?G             ]@�       �       
             �?�ȉo(��?9            �V@�       �                    X@�(\����?2             T@������������������������       �                     �?�       �                   �c@�Fǌ��?1            �S@�       �                   `a@������?             B@������������������������       �                     <@�       �                    �N@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                    �E@�       �                    �L@"pc�
�?             &@������������������������       �                      @�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �p@z�G�z�?             9@�       �                   @c@�q�q�?
             .@�       �                   l@      �?              @�       �                   �^@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     $@������������������������       �                     @�       �                    @K@^������?            �A@�       �                    �?j���� �?             1@������������������������       �                     @�       �                   �`@�q�q�?	             (@�       �                    �C@X�<ݚ�?             "@������������������������       �                     �?�       �                     F@      �?              @������������������������       �                     @�       �                    @���Q��?             @������������������������       �                      @�       �                   0k@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   0b@�����H�?             2@������������������������       �                     &@�       �                   ``@����X�?             @�       �                    �L@      �?             @������������������������       �                     �?�       �                   @_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?�Y闠��?o            �e@�       �                   �d@n�����?E            �\@�       �                   P`@X�;�^o�?B            �[@�       �       	          @33�? =[y��?,             Q@�       �                   0n@      �?              @�       �                    �?؇���X�?             @������������������������       �                     @�       �                   @\@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �? �.�?Ƞ?%             N@������������������������       �                     E@�       �                   s@�X�<ݺ?             2@������������������������       �                     1@������������������������       �                     �?�       �                   �b@0,Tg��?             E@������������������������       �                     *@�       �                    �?����"�?             =@�       �                   �i@��s����?             5@������������������������       �                      @�       �                   �d@�	j*D�?             *@�       �                    �?և���X�?             @�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?�       �                   �b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   `_@o����?*             M@�       �                    �P@���|���?             6@�       �                   @]@��
ц��?
             *@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       
             �?�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �       	          hff@tk~X��?             B@�       �                   �d@��hJ,�?             A@������������������������       �                     9@�       �       
             �?X�<ݚ�?             "@�       �                   �c@����X�?             @�       �       	          ����?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                      @ri  trj  bh�h"h#K �rk  h%�rl  Rrm  (KK�KK�rn  hV�B�        u@     �x@     �q@     �q@      *@     �W@      (@     �C@       @      �?              �?       @              $@      C@       @      ,@       @              @      ,@      @      ,@      �?      �?      �?                      �?       @      *@      �?      *@      �?      "@      �?      @              @      �?                      @              @      �?              @               @      8@      �?      2@              .@      �?      @      �?      �?              �?      �?                       @      �?      @              @      �?              �?      L@              F@      �?      (@              (@      �?             �p@      g@     �P@     @a@      I@      B@      8@      <@      8@      ,@      8@      &@      �?       @              �?      �?      @              @      �?              7@      @      @      @      @                      @      2@                      @              ,@      :@       @      9@      @      2@      @      @              &@      @              �?      &@      @              @      &@      �?      $@      �?              �?      $@              �?              @              �?      @              @      �?              1@     �Y@       @              .@     �Y@      @      "@      @              @      "@      �?       @      �?      @      �?                      @              @       @      �?              �?       @              "@     @W@      @      S@       @      *@              *@       @              @     �O@      �?      @              @      �?               @     �M@             �I@       @       @              @       @      @              @       @              @      1@      @      @       @               @      @              @       @                      (@      i@     �G@     �Q@      @      >@             �D@      @     �D@      @       @      �?       @                      �?     �C@      @     �B@      �?      *@              8@      �?      7@              �?      �?              �?      �?               @       @               @       @                      �?     @`@      E@     �]@      3@      &@      @      �?              $@      @      @      @      @      @      @              �?      @              @      �?                      @      @             �Z@      (@     �Z@      "@     �U@      @     �S@       @              �?     �S@      �?     �A@      �?      <@              @      �?      @                      �?     �E@              "@       @       @              �?       @               @      �?              4@      @      $@      @      @      @      @      �?              �?      @                      @      @              $@                      @      (@      7@      $@      @      @              @      @      @      @              �?      @      @      @               @      @               @       @      �?       @                      �?              @       @      0@              &@       @      @       @       @      �?              �?       @               @      �?                      @     �K@     �]@      2@     @X@      ,@      X@      @     @P@       @      @      �?      @              @      �?       @               @      �?              �?              �?     �M@              E@      �?      1@              1@      �?              &@      ?@              *@      &@      2@      @      1@               @      @      "@      @      @      @      �?              �?      @                       @              @      @      �?      @                      �?      @      �?      @                      �?     �B@      5@       @      ,@      @      @      @      �?      @                      �?              @      �?       @      �?                       @      =@      @      =@      @      9@              @      @       @      @       @       @       @                       @              @       @                       @ro  trp  bubhhubh)�rq  }rr  (hhh	h
hNhKhKhG        hh hNhJ	�tlhG        hNhG        h<Kh=Kh>h"h#K �rs  h%�rt  Rru  (KK�rv  hV�C              �?rw  trx  bhJhZhEC       ry  �rz  Rr{  h^Kh_h`Kh"h#K �r|  h%�r}  Rr~  (KK�r  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjMhkh"h#K �r�  h%�r�  Rr�  (KM�r�  hr�B�8         �                    �?�+	G�?�           ��@       g                    c@��4:���?�            Px@       @                   P`@ ˤ���?�            t@       %                    �?�Cc}h��?�             l@                          �Z@��
�π�?p            �d@                          �Z@؇���X�?!            �H@       
                   �Q@���}<S�?              G@       	                    �?      �?              @������������������������       �                     �?������������������������       �                     �?                          �\@t��ճC�?             F@                           �?      �?             @������������������������       �                      @������������������������       �                      @                           �?�(\����?             D@                           @G@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     A@������������������������       �                     @                           _@���#�İ?O            �]@                           `R@�Fǌ��?2            �S@������������������������       �        1            �S@������������������������       �                     �?       $                   �h@$�q-�?            �C@                          �_@���!pc�?	             &@              	          @33�?�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?      �?              @������������������������       �                     �?        !                    @H@؇���X�?             @������������������������       �                     @"       #                    @I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     <@&       /                   �_@F�t�K��?'            �L@'       .                   �Z@      �?              @(       )                    �?���Q��?             @������������������������       �                     �?*       +       	          ����?      �?             @������������������������       �                     �?,       -                    �O@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @0       ?                    �?�q��/��?!            �H@1       :                   �b@z�G�z�?             >@2       5       	             �?      �?             8@3       4                    _@      �?             @������������������������       �                      @������������������������       �                      @6       9                    �?P���Q�?             4@7       8                   0o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     2@;       <                    �L@      �?             @������������������������       �                      @=       >                    X@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     3@A       ^       
             �?R�L=��?:            @X@B       K                    @K@�ӭ�a��?,             R@C       D                   �a@`Jj��?             ?@������������������������       �                     *@E       J                   �b@�����H�?             2@F       I                   pb@����X�?             @G       H                    @E@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     &@L       U                   0i@��P���?            �D@M       P                    �?�eP*L��?             &@N       O                   �`@      �?             @������������������������       �                     �?������������������������       �                     @Q       T                   0f@����X�?             @R       S                   �b@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?V       Y       	          ����?ףp=
�?             >@W       X                    �?���Q��?             @������������������������       �                     @������������������������       �                      @Z       [                    @P@`2U0*��?             9@������������������������       �                     6@\       ]                   �k@�q�q�?             @������������������������       �                      @������������������������       �                     �?_       d                   0k@��H�}�?             9@`       a                    b@r�q��?
             2@������������������������       �                     ,@b       c                    �?      �?             @������������������������       �                     @������������������������       �                     �?e       f                    �L@؇���X�?             @������������������������       �                     @������������������������       �                     �?h       �                   `f@�������?'             Q@i       �                    @O@X�<ݚ�?&            �O@j       m                   j@|��?���?!             K@k       l                    �?r�q��?
             2@������������������������       �        	             .@������������������������       �                     @n       �                    �?<ݚ)�?             B@o       x                    �?r٣����?            �@@p       w                    b@      �?              @q       r                   �c@�q�q�?             @������������������������       �                     �?s       t                   �d@z�G�z�?             @������������������������       �                     @u       v       	          @33�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @y       ~                    b@�J�4�?             9@z       {                   �q@P���Q�?             4@������������������������       �                     0@|       }                    \@      �?             @������������������������       �                     �?������������������������       �                     @       �                   Pd@���Q��?             @������������������������       �                      @�       �                   `m@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     "@������������������������       �                     @�       �                    @L@bPD΂_�?�            �u@�       �       	          ����?��hJ,�?�            �m@�       �                    @G@���ۑ��?{            �h@�       �                   �c@��<b�ƥ?8             W@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �o@�E�����?6            �V@������������������������       �        &            �N@�       �                    �?XB���?             =@�       �                    �?���N8�?             5@������������������������       �                     @�       �                    �B@@4և���?             ,@�       �                     @@z�G�z�?             @������������������������       �                     @�       �                   @c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �                      @�       �                   �f@ ˤ���?C            �Z@�       �                    �G@(N:!���?B            @Z@�       �                   �_@�q�q�?             (@������������������������       �                      @�       �                   �]@z�G�z�?             $@������������������������       �                     �?�       �                   a@�����H�?             "@�       �                   �e@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    @��y� �?:            @W@�       �                   @Z@�X�<ݺ?9            �V@�       �                    �?�q�q�?             @�       �                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                   �Z@XB���?6            �U@�       �                   �X@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�D�e���?4            @U@������������������������       �                     G@�       �                     I@�7��?            �C@�       �                   �f@�<ݚ�?             "@������������������������       �                     �?�       �                   @p@      �?              @������������������������       �                     @�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     >@������������������������       �                     @������������������������       �                      @�       �                   �a@Hث3���?            �C@�       �                    �?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�       �       	             @��X��?             <@�       �                   `c@�㙢�c�?             7@�       �                    �?�����?             5@������������������������       �                     *@�       �                    �H@      �?              @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?n�tl��?C            �Z@�       �       	          ����?�i#[��?4             U@�       �                    �Q@�5��
J�?             G@�       �                   �T@�������?             F@������������������������       �                     �?�       �                    _@&^�)b�?            �E@�       �       
             �?և���X�?             @������������������������       �                     @�       �                     P@      �?             @������������������������       �                     @������������������������       �                     �?�       �       	          pff�?4?,R��?             B@�       �                   �a@ףp=
�?             >@������������������������       �                     3@�       �       	          ����?���!pc�?             &@�       �                    ^@      �?             @������������������������       �                      @�       �                   �m@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �a@�q�q�?             @������������������������       �                     @�       �                    @M@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �       
             �?���y4F�?             C@�       �                   @L@�X�<ݺ?	             2@������������������������       �                     �?������������������������       �                     1@�       �                    �Q@��Q��?             4@�       �                   0b@b�2�tk�?             2@�       �                    �?�8��8��?             (@�       �       	          `ff�?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    �?��<b���?             7@������������������������       �                     �?�                           @"pc�
�?             6@�       �                    �N@�KM�]�?             3@������������������������       �                     &@�       �                    �?      �?              @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       	             @z�G�z�?             @������������������������       �                     @������������������������       �                     �?            	          433�?�q�q�?             @������������������������       �                      @������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMKK�r�  hV�B0       `t@     �y@     �R@     �s@      E@     pq@      6@     @i@      &@     �c@      @      E@      @      E@      �?      �?              �?      �?              @     �D@       @       @       @                       @      �?     �C@      �?      @      �?                      @              A@      @              @     �\@      �?     �S@             �S@      �?              @      B@      @       @       @      �?              �?       @              �?      @              �?      �?      @              @      �?      �?      �?                      �?              <@      &@      G@      @      @       @      @              �?       @       @              �?       @      �?       @                      �?      @              @     �E@      @      8@      @      5@       @       @               @       @              �?      3@      �?      �?              �?      �?                      2@      @      @               @      @      �?      @                      �?              3@      4@     @S@      &@     �N@       @      =@              *@       @      0@       @      @      �?      @      �?                      @      �?                      &@      "@      @@      @      @      �?      @      �?                      @      @       @      @      �?      @                      �?              �?      @      ;@       @      @              @       @              �?      8@              6@      �?       @               @      �?              "@      0@      @      .@              ,@      @      �?      @                      �?      @      �?      @                      �?     �@@     �A@      <@     �A@      <@      :@      @      .@              .@      @              9@      &@      9@       @      @      @      @       @              �?      @      �?      @              �?      �?      �?                      �?               @      5@      @      3@      �?      0@              @      �?              �?      @               @      @               @       @      �?              �?       @                      @              "@      @             `o@     �W@     `i@     �A@     �f@      0@     �V@       @      �?      �?      �?                      �?     @V@      �?     �N@              <@      �?      4@      �?      @              *@      �?      @      �?      @              �?      �?              �?      �?              "@               @             @W@      ,@     @W@      (@       @      @               @       @       @              �?       @      �?       @      �?              �?       @              @             @U@       @     @U@      @      �?       @      �?      �?              �?      �?                      �?      U@      @      �?      �?      �?                      �?     �T@       @      G@             �B@       @      @       @              �?      @      �?      @              �?      �?      �?                      �?      >@                      @               @      4@      3@      �?      $@      �?                      $@      3@      "@      3@      @      3@       @      *@              @       @      @              �?       @               @      �?                       @              @      H@     �M@     �E@     �D@     �A@      &@     �A@      "@              �?     �A@       @      @      @      @              �?      @              @      �?              ?@      @      ;@      @      3@               @      @      @      @       @              �?      @              @      �?              @              @       @      @              �?       @      �?                       @               @       @      >@      �?      1@      �?                      1@      @      *@      @      &@      �?      &@      �?      @              @      �?                       @      @                       @      @      2@      �?              @      2@       @      1@              &@       @      @      �?       @      �?                       @      �?      @              @      �?               @      �?       @                      �?r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�ޡhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjMhkh"h#K �r�  h%�r�  Rr�  (KM�r�  hr�B�=         �                    @L@6������?�           ��@       M       	          ����?h�����?&            |@                          �Z@ά��.��?�            @p@                           �?����X�?	             ,@                           W@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @	                           �?"�W1��?�            �n@
                           @C@ �q�q�?.             R@                           �B@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?                          �`@�]0��<�?(            �N@                          ht@@3����?#             K@������������������������       �        !             I@                           @K@      �?             @������������������������       �                     �?������������������������       �                     @                          �`@؇���X�?             @                          @q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       "                   �c@�c�Α�?o            �e@       !                    b@      �?             6@                            �?D�n�3�?             3@                           @J@�8��8��?             (@������������������������       �                     @                           �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @#       ,                    �?�|�ʒ�?b             c@$       +                    @K@D�n�3�?             3@%       *                    �I@      �?             0@&       '                   Pc@�n_Y�K�?             *@������������������������       �                     @(       )                   i@z�G�z�?	             $@������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @-       B                    �?�������?T            �`@.       3                     E@��Zy�?            �C@/       2                    �B@z�G�z�?             $@0       1                    @A@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @4       A                    �?l��[B��?             =@5       >                    �?�û��|�?             7@6       =                   �t@p�ݯ��?             3@7       8                    @F@      �?
             0@������������������������       �                      @9       :                   �`@؇���X�?	             ,@������������������������       �                     &@;       <                    _@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @?       @                   `]@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @C       D                   �p@heu+��?;            �W@������������������������       �        .            �O@E       F                    @E@��a�n`�?             ?@������������������������       �                     .@G       L                    @     ��?             0@H       I                    �?"pc�
�?             &@������������������������       �                     @J       K                   �p@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @N       y                    �?V��N��?�            �g@O       P                    �F@�ص�ݒ�?U            @_@������������������������       �                     ?@Q       f       	          ����?t/*�?A            �W@R       _                    b@����"�?             =@S       T                    �?      �?             4@������������������������       �                     @U       ^                    @K@�t����?             1@V       ]                    �?      �?             0@W       X       	             �?$�q-�?	             *@������������������������       �                      @Y       \                    @G@�C��2(�?             &@Z       [                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?`       c                    �H@�q�q�?             "@a       b                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?d       e                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?g       n                    g@$�q-�?/            @P@h       i                   �U@     ��?
             0@������������������������       �                      @j       m                    �?@4և���?	             ,@k       l                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@o       p                   �m@@9G��?%            �H@������������������������       �                     6@q       v       
             �?�>����?             ;@r       u                    n@���7�?             6@s       t                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     4@w       x                    ]@z�G�z�?             @������������������������       �                     �?������������������������       �                     @z       �       	             @�9mf��?+            �O@{       �       
             �?��}*_��?%             K@|       �                    �?���!pc�?             F@}       ~                    �?@4և���?
             ,@������������������������       �                     &@       �                    c@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                     F@d��0u��?             >@������������������������       �                     @�       �                    @I@
;&����?             7@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     @�       �                   @^@������?             .@������������������������       �                     @�       �                    �?���|���?	             &@�       �                   0b@����X�?             @�       �                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �_@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �b@z�G�z�?             $@�       �                    �?�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     "@�       �                    �?��
n��?�            �q@�       �                   `]@��YIY�?m            �d@�       �                    �R@$Q�q�?,            �O@�       �                    �?�.ߴ#�?*            �N@�       �                    �L@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    x@���U�?&            �L@�       �                   0p@�h����?%             L@������������������������       �                     E@�       �                     P@@4և���?             ,@�       �                    �O@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       
             �?`Y�K�?A             Z@�       �                   pc@XB���?             =@������������������������       �                     2@�       �       	          ����?�C��2(�?             &@������������������������       �                     @�       �                    �N@r�q��?             @������������������������       �                     @�       �                   �t@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?�M;q��?.            �R@�       �                   �c@���|���?             6@�       �                    �?�z�G��?
             4@������������������������       �                     @�       �                   ``@      �?             0@�       �                     O@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   0d@"pc�
�?             &@������������������������       �                     @�       �                   �d@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    �?f1r��g�?#            �J@�       �                    ^@������?             A@�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   �a@z�G�z�?             @������������������������       �                      @�       �                    @N@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       
             �?؇���X�?             <@�       �                    @N@      �?             0@�       �                   b@���Q��?             @�       �                   �[@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   �h@�C��2(�?             &@�       �                   �R@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �                     (@������������������������       �                     3@�       �                   �^@���k��?M            �]@�       �                    �?������?            �D@�       �                    �?���Q��?             >@�       �       	             �?�z�G��?             $@������������������������       �                     @�       �                   `X@���Q��?             @������������������������       �                      @�       �                   �u@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                     N@      �?             4@�       �                    @M@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   `a@�r����?             .@�       �                    @R@����X�?             @�       �                    k@r�q��?             @������������������������       �                     @�       �                   Po@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     &@�       �                   `Q@���L��?2            �S@�       �                   �`@r�q��?             (@�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@�       �                   �f@�X����?,            �P@������������������������       �                     @�             	          ����?:���W�?(            �M@�             
             �?���N8�?             E@�                         �c@z�G�z�?             D@�       �                   �a@�>����?             ;@������������������������       �        	             (@                         �a@�r����?
             .@������������������������       �                     �?            	            �?@4և���?	             ,@                         `@r�q��?             @                        �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @	                        `d@��
ц��?	             *@
                         �P@      �?              @                        �]@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                        `]@ҳ�wY;�?             1@            	          hff @      �?             @������������������������       �                     @������������������������       �                     �?                        �l@�θ�?	             *@            	          pff�?���Q��?             @������������������������       �                     �?            	          033@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMKK�r�  hV�B�       �t@     �x@      o@     �h@     �h@     �N@      @      $@      @      @              @      @                      @     `h@     �I@     @Q@      @      $@      �?      $@                      �?     �M@       @     �J@      �?      I@              @      �?              �?      @              @      �?      �?      �?              �?      �?              @             �_@      H@      &@      &@      &@       @      &@      �?      @              @      �?      @                      �?              @              @     �\@     �B@      &@       @       @       @       @      @              @       @       @               @       @                      @      @              Z@      =@      1@      6@       @       @       @      �?              �?       @                      @      .@      ,@      "@      ,@      @      (@      @      (@       @               @      (@              &@       @      �?              �?       @              @               @       @               @       @              @             �U@      @     �O@              8@      @      .@              "@      @      "@       @      @              @       @               @      @                      @      I@     @a@      0@     @[@              ?@      0@     �S@      &@      2@      @      .@      @               @      .@      �?      .@      �?      (@               @      �?      $@      �?       @               @      �?                       @              @      �?              @      @      @      �?      @                      �?      �?       @               @      �?              @      N@      @      *@       @              �?      *@      �?       @               @      �?                      &@       @     �G@              6@       @      9@      �?      5@      �?      �?              �?      �?                      4@      �?      @      �?                      @      A@      =@      A@      4@      @@      (@      *@      �?      &@               @      �?              �?       @              3@      &@      @              (@      &@      �?      @      �?                      @      &@      @      @              @      @      @       @      �?       @               @      �?              @               @       @               @       @               @       @      �?       @      �?                       @      �?                      "@     �U@      i@      ;@     �a@      @     �M@      @      M@      �?      @      �?                      @       @     �K@      �?     �K@              E@      �?      *@      �?      @              @      �?                      "@      �?              �?      �?      �?                      �?      7@     @T@      �?      <@              2@      �?      $@              @      �?      @              @      �?      �?              �?      �?              6@     �J@      ,@       @      ,@      @      @              $@      @      �?      @              @      �?              "@       @      @              @       @               @      @                       @       @     �F@       @      :@      @       @              �?      @      �?       @               @      �?              �?       @              @      8@      @      (@      @       @      �?       @      �?                       @       @              �?      $@      �?      �?              �?      �?                      "@              (@              3@     �M@      N@      (@      =@      (@      2@      @      @      @               @      @               @       @      �?       @                      �?      @      .@      @       @               @      @               @      *@       @      @      �?      @              @      �?      �?      �?                      �?      �?                       @              &@     �G@      ?@       @      $@       @      �?       @                      �?              "@     �F@      5@      @              C@      5@      @@      $@      @@       @      9@       @      (@              *@       @              �?      *@      �?      @      �?      �?      �?      �?                      �?      @               @              @      @       @      @      �?      @      �?                      @      �?              @                       @      @      &@      @      �?      @                      �?      @      $@      @       @              �?      @      �?      @                      �?               @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJQY%hG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjMhkh"h#K �r�  h%�r�  Rr�  (KM�r�  hr�B�9         �       	          ����?�Z���?�           ��@       G                    �?�q�q�?�             x@              	          `ffֿ���ѽ��?`             d@������������������������       �                     @                           @D@���@M^�?[            `c@������������������������       �        
             3@                           �?�ʻ����?Q             a@                          �a@�<ݚ�?             ;@	       
                   �`@���Q��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     1@       <                    �?\��bi�?E            @[@       '                   �`@7�A�0�?7             V@                            a@ҐϿ<��?'            �N@                           �?tk~X��?             B@                          �_@$�q-�?             :@������������������������       �                     (@                           �?؇���X�?             ,@������������������������       �                     �?                           `@8�Z$���?             *@                            I@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @                           @P@      �?             $@                           Z@����X�?             @                           \@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @!       "                   Pb@� �	��?             9@������������������������       �                     (@#       $                   �c@8�Z$���?
             *@������������������������       �                     @%       &                   �n@�q�q�?             @������������������������       �                      @������������������������       �                     @(       -                   �d@�5��?             ;@)       *                    T@      �?              @������������������������       �                     @+       ,                    �?      �?             @������������������������       �                     @������������������������       �                     �?.       7                    k@���y4F�?             3@/       6       	          @33�?և���X�?             @0       5                     N@      �?             @1       2                     K@      �?             @������������������������       �                     �?3       4                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?8       ;                    �I@�8��8��?             (@9       :                    �G@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @=       B       	          ����?�����?             5@>       ?                   �^@�X�<ݺ?             2@������������������������       �                     $@@       A                    �G@      �?              @������������������������       �                     �?������������������������       �                     @C       F       
             �?�q�q�?             @D       E                    ]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?H       U                    @G@�1c�#�?�            �k@I       P                    @x�G�z�?4             T@J       O                    �A@�"w����?1             S@K       N                   �\@$�q-�?
             *@L       M                    �@@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �        '            �O@Q       R       
             �?      �?             @������������������������       �                     �?S       T                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?V       [                   �\@�o{�88�?^            �a@W       X                   �j@���|���?	             &@������������������������       �                     @Y       Z                   �m@z�G�z�?             @������������������������       �                     @������������������������       �                     �?\       a                    I@\|/��j�?U            �`@]       ^                    �?���Q��?             $@������������������������       �                      @_       `                    �?      �?              @������������������������       �                     @������������������������       �                     @b       c                   @k@��̋���?O            �^@������������������������       �                     B@d       �                    �?�4���L�?5            �U@e       ~                    @     ��?1             T@f       }                   `g@�J�4�?.            �R@g       l                    �?�x
�2�?-            �R@h       k                   0b@���N8�?             5@i       j                    @O@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             .@m       v       	            �?r�����?             �J@n       o                   pa@������?            �D@������������������������       �                     $@p       u                    @I@��� ��?             ?@q       r                   �^@և���X�?             @������������������������       �                      @s       t                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     8@w       |                   xp@      �?             (@x       y                    _@      �?              @������������������������       �                     @z       {                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?       �                    �N@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    `@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    �?��E�V�?�            �u@�       �                    �?���k�6�?�            @o@�       �                    `P@�v:���?(             Q@�       �                   �c@Nd^����?$            �N@�       �                    �?�`���?            �H@�       �                   �a@ҳ�wY;�?             A@�       �                   �`@      �?             6@�       �                    @H@"pc�
�?             &@������������������������       �                     �?�       �                    �J@ףp=
�?             $@������������������������       �                      @�       �                    `@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   @b@"pc�
�?             &@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @�       �       	             �?      �?             @������������������������       �                      @������������������������       �                      @�       �                   pc@�8��8��?	             (@������������������������       �                     $@�       �                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          `ff�?z�G�z�?
             .@�       �                    �?և���X�?             @�       �                   @]@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@������������������������       �                     @�       �                    @G@d}h���?~            �f@�       �                   �`@b�2�tk�?             B@������������������������       �        	             0@�       �                   (p@�z�G��?             4@�       �                   �b@@�0�!��?             1@�       �                   Pm@���!pc�?             &@�       �                    �?      �?             @������������������������       �                      @�       �                   �\@      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   �i@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    @J@��-*�?h            @b@�       �                   @c@ 7���B�?             ;@������������������������       �                     7@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �J@J��ԛ�?T            �]@�       �       
             �?�q�q�?             "@������������������������       �                     �?�       �       	          ����?      �?              @������������������������       �                      @�       �                    c@�q�q�?             @�       �                    �?z�G�z�?             @�       �                   p`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                   �_@�2����?N            �[@�       �                   @_@�����?-            �P@�       �                   �s@(;L]n�?)             N@�       �                   `X@ _�@�Y�?'             M@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �        !             I@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                   �h@8�$�>�?!            �E@�       �                    �K@      �?              @������������������������       �                     �?�       �                   0`@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                   pb@��R[s�?            �A@�       �                   �p@     ��?             @@�       �                    �L@�}�+r��?             3@�       �                   �d@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@�       �                    �?�n_Y�K�?             *@������������������������       �                     @�       �                   �\@����X�?             @������������������������       �                     �?�       �                    �?r�q��?             @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �? "��u�?C             Y@�       �                    �?      �?              @������������������������       �                     @�       �                    �N@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    `@�nkK�?=             W@������������������������       �                     <@�                          @s@      �?(             P@�       �                   �b@h�����?#             L@������������������������       �        !            �J@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                         �P@      �?              @                         �L@؇���X�?             @������������������������       �                     @                         �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMKK�r�  hV�Bp        u@     �x@     @o@     �`@      N@     @Y@              @      N@     �W@              3@      N@      S@      5@      @      @      @      @                      @      1@             �C@     �Q@     �B@     �I@      5@      D@      @      =@       @      8@              (@       @      (@              �?       @      &@       @      @              @       @                      @      @      @      @       @      �?       @      �?                       @      @                      @      ,@      &@      (@               @      &@              @       @      @       @                      @      0@      &@      �?      @              @      �?      @              @      �?              .@      @      @      @      @      @      @      �?      �?               @      �?       @                      �?               @      �?              &@      �?      @      �?      @                      �?       @               @      3@      �?      1@              $@      �?      @      �?                      @      �?       @      �?      �?              �?      �?                      �?     �g@     �@@     @S@      @     �R@      �?      (@      �?      �?      �?      �?                      �?      &@             �O@               @       @              �?       @      �?       @                      �?     @\@      >@      @      @              @      @      �?      @                      �?     @[@      7@      @      @               @      @      @      @                      @     @Z@      1@      B@             @Q@      1@     @P@      .@     �O@      (@     �O@      &@      4@      �?      @      �?              �?      @              .@             �E@      $@     �B@      @      $@              ;@      @      @      @               @      @       @               @      @              8@              @      @       @      @              @       @       @       @                       @      @                      �?       @      @              @       @              @       @               @      @              V@     `p@     �T@      e@     �E@      9@      B@      9@      8@      9@      (@      6@      &@      &@      "@       @              �?      "@      �?       @              �?      �?              �?      �?               @      "@              @       @      @               @       @       @       @                       @      �?      &@              $@      �?      �?              �?      �?              (@      @      @      @      @      �?              �?      @              �?       @               @      �?               @              (@              @             �C@     �a@      ,@      6@              0@      ,@      @      ,@      @       @      @      @      @       @              �?      @              �?      �?       @              �?      �?      �?      �?                      �?      @              @                      @      9@     @^@      �?      :@              7@      �?      @              @      �?              8@     �W@      @      @              �?      @       @       @              @       @      @      �?       @      �?              �?       @               @                      �?      2@      W@      @      P@       @      M@      �?     �L@      �?      @              @      �?                      I@      �?      �?              �?      �?              �?      @      �?                      @      .@      <@      @       @              �?      @      �?              �?      @              "@      :@      @      :@      �?      2@      �?      @              @      �?                      .@      @       @              @      @       @              �?      @      �?      �?      �?              �?      �?              @              @              @     �W@       @      @              @       @      �?       @                      �?      @      V@              <@      @      N@       @      K@             �J@       @      �?              �?       @               @      @      �?      @              @      �?      @      �?                      @      �?        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ��fbhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjK�hkh"h#K �r�  h%�r�  Rr�  (KK�r�  hr�BH4         �                    �?�#i����?�           ��@       M       	          ����?D�X%��?           �x@                          �_@� e��?[            �a@              
             �?�L���?            �B@                          �_@      �?             @@������������������������       �                     4@                           �I@�8��8��?
             (@       	                    �?r�q��?             @������������������������       �                     �?
                           �?z�G�z�?             @                          a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @                          �_@���Q��?             @������������������������       �                      @                           �M@�q�q�?             @������������������������       �                     �?������������������������       �                      @       $                    �?^%�e��?A            �Z@                           �F@��
ц��?             :@������������������������       �                     @                           �?և���X�?             5@������������������������       �                     @       #                    �N@X�Cc�?
             ,@       "                    @M@      �?             $@       !       	             �?X�<ݚ�?             "@                           Z@      �?              @������������������������       �                      @                           Pf@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @%       6                   �b@     ��?0             T@&       5                   �p@�q�q��?             H@'       4       	          ����?p9W��S�?             C@(       1                   �_@�G��l��?             5@)       .                   p`@z�G�z�?             $@*       +                    �?      �?              @������������������������       �                     @,       -                   �k@�q�q�?             @������������������������       �                     �?������������������������       �                      @/       0                   0a@      �?              @������������������������       �                     �?������������������������       �                     �?2       3                    �J@���!pc�?             &@������������������������       �                      @������������������������       �                     @������������������������       �                     1@������������������������       �                     $@7       >                   �^@     ��?             @@8       9                   pi@�z�G��?             $@������������������������       �                     @:       =                    e@      �?             @;       <                   pc@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @?       F                   �a@�X����?             6@@       E                   Pd@�8��8��?             (@A       D       	             �?      �?             @B       C                     L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @G       H                   �f@���Q��?             $@������������������������       �                     @I       J                   �b@؇���X�?             @������������������������       �                     @K       L                     E@      �?              @������������������������       �                     �?������������������������       �                     �?N       O                   �U@�m(�X�?�            �o@������������������������       �                     �?P                           �?HVĮ���?�            �o@Q       v       	          pff�?l������?v             e@R       q                   pc@�Y�����?8            �T@S       n       	          ����?z���=��?4            @S@T       _                    �?d1<+�C�?2            @R@U       V                   `_@�IєX�?$            �I@������������������������       �                     8@W       Z                   �[@�����H�?             ;@X       Y       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @[       ^                    @H@ �q�q�?             8@\       ]                    �E@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     5@`       m                   �_@�X����?             6@a       l                    ^@���y4F�?             3@b       i       	          033�?����X�?             ,@c       d                    @K@      �?             @������������������������       �                      @e       f                    �?      �?             @������������������������       �                      @g       h                   �X@      �?              @������������������������       �                     �?������������������������       �                     �?j       k                    �N@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @o       p                    �?      �?             @������������������������       �                     @������������������������       �                     �?r       s                   �d@�q�q�?             @������������������������       �                     @t       u                    b@�q�q�?             @������������������������       �                      @������������������������       �                     �?w       ~       	          `ff @�D�e���?>            @U@x       }                   �d@@-�_ .�?            �B@y       z                    @J@      �?             @������������������������       �                     �?{       |                   �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                    �@@������������������������       �        !             H@�       �                    Y@��f�{��?1            �U@�       �                    �?�����H�?             "@�       �                    k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        +            @S@�       �                    �?,Tg�x0�?�             u@�       �                   `c@�̐d��?>            @Z@�       �                   �Q@ p�/��?7            @V@������������������������       �                     �?�       �                   �Z@�zvܰ?6             V@�       �                   �X@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �n@�D�e���?3            @U@������������������������       �                    �I@�       �                    o@�IєX�?             A@������������������������       �                     �?�       �                    @I@Pa�	�?            �@@�       �                   �q@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     <@�       �                    �?     ��?             0@�       �                   v@      �?              @������������������������       �                     @������������������������       �                      @�       �                   �]@      �?              @������������������������       �                     �?������������������������       �                     @�       �                    Z@��cv�?�            �l@������������������������       �                     @�       �                    @L@���x��?�            @l@�       �       	          ����?�E���-�?[             b@�       �       	          ����?@-�_ .�?E            �[@�       �                    I@����?A            �Z@�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   Pr@ ��WV�??             Z@�       �                    @p�C��?9            �V@�       �                   @[@�E�����?8            �V@�       �                    ]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        6             V@������������������������       �                     �?�       �                    @8�Z$���?             *@������������������������       �                     &@������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �d@�'�=z��?            �@@������������������������       �                     @�       �       
             �?�n_Y�K�?             :@������������������������       �                     @�       �                     F@      �?             4@�       �       	             @؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    �K@�	j*D�?             *@�       �                    �?�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �       
             �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �_@D^��#��?4            �T@�       �                    �?�z�G��?             4@������������������������       �                     @�       �                    �?���Q��?             .@�       �                    �M@r�q��?             @�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �       	          ����?�g�y��?%             O@�       �                   �O@¦	^_�?             ?@������������������������       �                     @�       �       	          ����?�+$�jP�?             ;@�       �                   �a@����X�?	             ,@�       �                    �?      �?             @�       �                    b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   Pc@ףp=
�?             $@������������������������       �                      @�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �q@$�q-�?	             *@������������������������       �                     &@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   pb@�4�����?             ?@�       �                   P`@�KM�]�?             3@������������������������       �                      @������������������������       �        
             1@�       �                    �?�q�q�?             (@�       �                   @\@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hV�B�       `u@     �x@     �V@     0s@     �Q@     @R@      @      A@      �?      ?@              4@      �?      &@      �?      @              �?      �?      @      �?       @      �?                       @               @              @       @      @               @       @      �?              �?       @             �P@     �C@      (@      ,@              @      (@      "@      @              @      "@      @      @      @      @      @      @       @               @      @              @       @                      �?      �?                      @     �K@      9@     �B@      &@      ;@      &@      $@      &@       @       @      �?      @              @      �?       @      �?                       @      �?      �?      �?                      �?       @      @       @                      @      1@              $@              2@      ,@      @      @              @      @      @      @      �?              �?      @                       @      .@      @      &@      �?      @      �?      �?      �?      �?                      �?       @               @              @      @      @              �?      @              @      �?      �?              �?      �?              5@     @m@      �?              4@     @m@      3@     �b@      1@     �P@      *@      P@      $@     �O@      @      H@              8@      @      8@       @      �?              �?       @              �?      7@      �?       @               @      �?                      5@      @      .@      @      .@      @      $@      @      @               @      @      �?       @              �?      �?      �?                      �?      �?      @              @      �?                      @      @              @      �?      @                      �?      @       @      @              �?       @               @      �?               @     �T@       @     �A@       @       @      �?              �?       @               @      �?                     �@@              H@      �?     @U@      �?       @      �?      �?              �?      �?                      @             @S@     `o@     @U@      W@      *@     @U@      @              �?     @U@      @       @      �?       @                      �?     �T@       @     �I@              @@       @              �?      @@      �?      @      �?      @                      �?      <@              @      "@      @       @      @                       @      �?      @      �?                      @     �c@      R@              @     �c@     �P@     @^@      7@     @Z@      @     @Y@      @      �?      �?              �?      �?              Y@      @     @V@       @     @V@      �?      �?      �?      �?                      �?      V@                      �?      &@       @      &@                       @      @      �?      @                      �?      0@      1@              @      0@      $@      @              $@      $@      @      �?      @                      �?      @      "@      �?       @               @      �?              @      �?      @                      �?      C@      F@      @      ,@              @      @      "@      @      �?      �?      �?      �?                      �?      @              �?       @               @      �?              @@      >@      6@      "@              @      6@      @      $@      @      �?      @      �?      �?      �?                      �?               @      "@      �?       @              �?      �?              �?      �?              (@      �?      &@              �?      �?              �?      �?              $@      5@       @      1@       @                      1@       @      @      @      �?              �?      @               @      @              @       @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ$�phG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r   tr  bK�r  Rr  }r  (hKhjK�hkh"h#K �r  h%�r  Rr  (KK�r  hr�B�2         �                    �?"��G,�?�           ��@       -                    �?Z�����?Y           ��@                           @K@|�-蝉�?W            �`@                           �?���!���?6            �S@                          `c@�LQ�1	�?             7@                           �G@      �?             4@                          �b@�q�q�?             @������������������������       �                     @	       
                    �?�q�q�?             @������������������������       �                     �?                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                          �Z@@4և���?             ,@������������������������       �                     �?������������������������       �                     *@������������������������       �                     @                          �q@�h����?'             L@������������������������       �                      F@                           �?�8��8��?             (@������������������������       �                     @                          �r@      �?              @������������������������       �                     �?������������������������       �                     @       &                    �?l��
I��?!             K@       #                    �?�X����?             6@       "                     Q@�z�G��?             4@                          ``@�<ݚ�?             2@������������������������       �                     @       !                   �a@��S�ۿ?	             .@                            �M@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �                      @$       %                    `@      �?              @������������������������       �                     �?������������������������       �                     �?'       (                    �?      �?             @@������������������������       �                     (@)       *       	          pff�?P���Q�?             4@������������������������       �        	             .@+       ,       	             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @.       E                    _@�Qrc_�?           p{@/       0                   `\@@�r-��?#            �M@������������������������       �        
             1@1       >                    �?d}h���?             E@2       3                    �?8����?             7@������������������������       �                     @4       =                    �?b�2�tk�?             2@5       :                    �?8�Z$���?	             *@6       7                   `@؇���X�?             @������������������������       �                     @8       9                   @M@�q�q�?             @������������������������       �                     �?������������������������       �                      @;       <                   @b@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @?       B       	          433�?�KM�]�?             3@@       A                    �O@�q�q�?             @������������������������       �                      @������������������������       �                     �?C       D                    ]@      �?	             0@������������������������       �                     �?������������������������       �                     .@F       �       	             �?0��'A�?�            �w@G       b                    �? �2�^�?p            �g@H       a                   �f@X3_��?(            �Q@I       V                   �b@�ՙ/�?%            �O@J       K       
             �?�xGZ���?            �A@������������������������       �                     @L       U       
             �?J�8���?             =@M       T       	          ����?\X��t�?             7@N       O                   �_@�q�q�?
             .@������������������������       �                     "@P       S                   0a@r�q��?             @Q       R                    @G@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @W       Z                   �`@�>4և��?             <@X       Y                    �B@�X�<ݺ?	             2@������������������������       �                     �?������������������������       �                     1@[       \                   �c@���Q��?             $@������������������������       �                      @]       ^                   �d@      �?              @������������������������       �                     @_       `                   l@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @c       j                   �_@�Y>J��?H            @]@d       g                   @]@8^s]e�?             =@e       f                     N@      �?             0@������������������������       �                     .@������������������������       �                     �?h       i                    b@�n_Y�K�?             *@������������������������       �                     @������������������������       �                      @k       v                   `]@��|���?;             V@l       m       
             �?X�<ݚ�?             "@������������������������       �                     �?n       o                   `b@      �?              @������������������������       �                     �?p       q                    �?����X�?             @������������������������       �                     �?r       s                    c@r�q��?             @������������������������       �                     @t       u                   �d@�q�q�?             @������������������������       �                     �?������������������������       �                      @w       �                   �t@$��$�L�?5            �S@x       �                    f@�:�^���?4            �S@y       |                   �c@�S(��d�?3            @S@z       {                    �?      �?              @������������������������       �                     �?������������������������       �                     �?}       �       	            �?��S�ۿ?1            �R@~                           �? ������?*            �O@������������������������       �        %            �L@�       �                    @L@r�q��?             @������������������������       �                     @�       �                   �g@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    _@�q�q�?             (@������������������������       �                      @�       �                   Pn@z�G�z�?             $@�       �                    �L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �       	          033�?r�q��?o             h@�       �                     F@�	j*D�?8            �V@�       �                    �?      �?              @�       �                    �D@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   `_@U7W1�?2            �T@������������������������       �                     C@�       �                    �?��S���?            �F@�       �                   �i@������?             >@������������������������       �                     @�       �                   pv@H%u��?             9@�       �       	          ����?�nkK�?             7@�       �                   a@�8��8��?             (@������������������������       �                     $@�       �                    �K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �                      @�       �                    �K@�r����?	             .@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@�       �                   pe@(a��䛼?7            @Y@�       �                   Pe@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �                    �?�nkK�?2             W@�       �       
             �?      �?&             P@�       �                    [@ ��WV�?             :@������������������������       �                     �?������������������������       �                     9@�       �                    @M@P�Lt�<�?             C@������������������������       �                    �@@�       �                     N@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �_@@4և���?             <@�       �                    p@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �        
             7@�       �       
             �?�+$�jP�?e            @d@�       �                    �J@$��m��?             :@������������������������       �                     @�       �                    �?��+7��?             7@������������������������       �                     (@�       �                   �a@�eP*L��?             &@�       �       	          ���ٿr�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    b@z�G�z�?             @������������������������       �                     @�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?��>z��?W             a@�       �                    y@��s��?=            �W@�       �                   ``@��<b�ƥ?;             W@������������������������       �        "            �H@�       �       	          ����? �#�Ѵ�?            �E@�       �                   �b@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     C@�       �                     L@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?v�2t5�?            �D@�       �       	             �?�G��l��?             5@�       �                   �\@      �?	             (@������������������������       �                     �?�       �                   0j@"pc�
�?             &@������������������������       �                      @������������������������       �                     "@�       �                    \@�����H�?             "@������������������������       �                     @�       �                    o@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �l@��Q��?             4@�       �                   p`@j���� �?             1@������������������������       �                     @�       �       	            �?r�q��?             (@�       �                   �h@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@������������������������       �                     @r	  tr
  bh�h"h#K �r  h%�r  Rr  (KK�KK�r  hV�B�       @s@     �z@     `q@     `r@      [@      9@     �Q@      "@      .@       @      .@      @       @      @              @       @      �?      �?              �?      �?              �?      �?              *@      �?              �?      *@                      @     �K@      �?      F@              &@      �?      @              @      �?              �?      @              C@      0@      @      .@      @      ,@      @      ,@      @              �?      ,@      �?      @              @      �?                      &@       @              �?      �?              �?      �?              ?@      �?      (@              3@      �?      .@              @      �?              �?      @             @e@     �p@      "@      I@              1@      "@     �@@      @      0@              @      @      &@       @      &@      �?      @              @      �?       @      �?                       @      �?      @              @      �?              @               @      1@      �?       @               @      �?              �?      .@      �?                      .@      d@     `k@     �_@     �N@      @@     �C@      8@     �C@      3@      0@              @      3@      $@      *@      $@      @      $@              "@      @      �?       @      �?              �?       @              @               @              @              @      7@      �?      1@      �?                      1@      @      @       @               @      @              @       @       @               @       @               @             �W@      6@      4@      "@      .@      �?      .@                      �?      @       @      @                       @     �R@      *@      @      @      �?              @      @      �?               @      @      �?              �?      @              @      �?       @      �?                       @     �Q@       @     �Q@      @     �Q@      @      �?      �?      �?                      �?     �Q@      @      O@      �?     �L@              @      �?      @              �?      �?      �?                      �?       @      @               @       @       @      �?       @               @      �?              @                      �?              �?      A@     �c@      <@     �O@      @      �?       @      �?              �?       @              @              5@      O@              C@      5@      8@       @      6@      @              @      6@      �?      6@      �?      &@              $@      �?      �?      �?                      �?              &@       @              *@       @      �?       @      �?                       @      (@              @     �W@       @      @              @       @              @      V@       @      O@      �?      9@      �?                      9@      �?     �B@             �@@      �?      @      �?                      @       @      :@       @      @              @       @                      7@      >@     �`@      "@      1@      @              @      1@              (@      @      @      @      �?              �?      @              �?      @              @      �?      �?      �?                      �?      5@     �\@      @     �V@       @     �V@             �H@       @     �D@       @      @       @                      @              C@       @      �?              �?       @              1@      8@      $@      &@      "@      @              �?      "@       @               @      "@              �?       @              @      �?      @      �?                      @      @      *@      @      $@      @               @      $@       @      �?       @                      �?              "@              @r  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJW:+LhG        hNhG        h<Kh=Kh>h"h#K �r  h%�r  Rr  (KK�r  hV�C              �?r  tr  bhJhZhEC       r  �r  Rr  h^Kh_h`Kh"h#K �r  h%�r  Rr  (KK�r  hE�C       r   tr!  bK�r"  Rr#  }r$  (hKhjMhkh"h#K �r%  h%�r&  Rr'  (KM�r(  hr�Bh:         f                   �`@�#i����?�           ��@       M                    �?p�L���?�            `s@       $       	          ����?H0sE�d�?�             l@              
             �?R�}e�.�?%             J@                          �Z@>A�F<�?             C@              	             пX�<ݚ�?             "@������������������������       �                     �?              	          hff�?      �?              @	       
                    @L@և���X�?             @������������������������       �                      @                          �[@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?                          �`@ܷ��?��?             =@������������������������       �                     1@                           _@      �?             (@                           \@ףp=
�?             $@                          �\@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                          @V@      �?
             ,@������������������������       �                     @                           �H@�z�G��?	             $@������������������������       �                     �?       #                    �?�<ݚ�?             "@                          @_@����X�?             @������������������������       �                     @       "                    �P@      �?             @        !                    [@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @%       :                    �?���y�?p            �e@&       7                   �z@�94�s0�?N            �\@'       6                   �^@ T���v�?L            @\@(       )                   @Z@l��\��?             A@������������������������       �                      @*       5                   Hs@ȵHPS!�?             :@+       .                    �?HP�s��?             9@,       -                   �l@�q�q�?             @������������������������       �                      @������������������������       �                     �?/       0                   `_@���7�?             6@������������������������       �                     2@1       4       	              @      �?             @2       3                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �        2            �S@8       9                   ��@      �?              @������������������������       �                     �?������������������������       �                     �?;       J                   P`@ܷ��?��?"             M@<       I                   �`@�NW���?             �J@=       H                   `^@z�G�z�?             4@>       ?                    �?      �?              @������������������������       �                      @@       G                   �p@�q�q�?             @A       B                   �Y@      �?             @������������������������       �                     �?C       D                   �j@�q�q�?             @������������������������       �                     �?E       F                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     (@������������������������       �                    �@@K       L                   �`@���Q��?             @������������������������       �                     @������������������������       �                      @N       a       	          ����?k�q��?7            @U@O       T                   `T@���Q��?&             N@P       S                    �?�z�G��?             4@Q       R                    \@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             *@U       ^                    �?      �?             D@V       W                    �L@z�G�z�?            �A@������������������������       �                     5@X       ]                   �o@      �?             ,@Y       \                   �j@�<ݚ�?             "@Z       [                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @_       `                     J@���Q��?             @������������������������       �                      @������������������������       �                     @b       c                     P@H%u��?             9@������������������������       �                     0@d       e                    �?�q�q�?             "@������������������������       �                     @������������������������       �                     @g       �                    �L@������?
           �z@h       �                    �?z�G��?�             t@i       j                   �G@��+-l�?�            �q@������������������������       �                      @k       �                    �?T�iA�?�            �q@l       �                    @L@@�&b
}�?4            �U@m       r                   �e@�Q����?1             T@n       o                   @[@z�G�z�?             $@������������������������       �                     �?p       q                    @K@�����H�?             "@������������������������       �                      @������������������������       �                     �?s       �                    �?և���X�?+            �Q@t       u                    @C@N1���?&            �N@������������������������       �                     @v       �                   `c@>4և���?#             L@w       �       	          ����?b�2�tk�?!             K@x       �                   8|@      �?             B@y       ~                   �o@4�2%ޑ�?            �A@z       }                   �h@�8��8��?	             (@{       |                    @J@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@       �                    `@8����?             7@�       �                    �J@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �?@�0�!��?             1@�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �p@�r����?             .@������������������������       �                      @������������������������       �                     *@������������������������       �                     �?�       �                    �F@�q�q�?             2@�       �                   pc@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �       
             �?8�Z$���?             *@������������������������       �                     @�       �                    �?      �?              @�       �                   Pn@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �l@z�G�z�?             @������������������������       �                     @�       �                    �J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �I@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?�ը
q��?{             h@������������������������       �                     ;@�       �                    @4�{Y���?h            �d@�       �       	             @��2(&�?`            @c@�       �                    �?�����?\            `b@�       �                    �?Ћ����?4            �T@�       �                   `o@0z�(>��?-            �Q@������������������������       �                    �E@�       �                    �B@ �Cc}�?             <@�       �                   @c@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   @_@`2U0*��?             9@�       �                   `p@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �        
             0@������������������������       �                     &@�       �       	          033�?�z����?(            @P@�       �                   `a@��� ��?&             O@�       �                   `]@��<D�m�?            �H@�       �                    @H@R���Q�?             4@�       �                   @[@��S�ۿ?             .@�       �                    �F@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@�       �                   �d@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     =@�       �                    �I@�n_Y�K�?             *@�       �                   �d@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?�q�q�?             (@������������������������       �                      @�       �       	          `ff�?�z�G��?             $@������������������������       �                     @�       �       
             �?      �?             @�       �                    �C@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �G@�s��:��?             C@������������������������       �                     "@�       �                   �c@�f7�z�?             =@�       �       	          ����?X�Cc�?	             ,@�       �                   �r@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �       	          `ffֿz�G�z�?             .@������������������������       �                     �?�       �                   �O@؇���X�?             ,@������������������������       �                      @������������������������       �                     (@�       �                   �_@��
ц��?D             Z@�       �                    �?     ��?             @@�       �                   c@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?             <@������������������������       �                     ,@�       �                   `Z@      �?
             ,@������������������������       �                     @�       �                    �?���|���?             &@�       �       	          033@�z�G��?             $@�       �                   �p@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�                         �c@)O���?.             R@�       �                    �?X�Emq�?!            �J@�       �       
             �?X�<ݚ�?            �F@�       �                     P@~�4_�g�?             F@�       �                   �a@����X�?            �A@�       �                   0q@��.k���?
             1@�       �       	          `ff�?�z�G��?             $@�       �                    @O@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �c@����X�?             @������������������������       �                     @������������������������       �                      @�       �                    �O@�����H�?             2@������������������������       �                     *@�       �                   `b@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     "@������������������������       �                     �?             	          ����?      �?              @������������������������       �                     @������������������������       �                     @                         r@���y4F�?             3@                         b@��S�ۿ?
             .@������������������������       �                     *@            
             �?      �?              @������������������������       �                     �?������������������������       �                     �?	      
                   �?      �?             @������������������������       �                     @������������������������       �                     �?r)  tr*  bh�h"h#K �r+  h%�r,  Rr-  (KMKK�r.  hV�B�       `u@     �x@     �O@     �n@      8@      i@      ,@      C@      @      ?@      @      @              �?      @      @      @      @               @      @      �?              �?      @                      �?      @      :@              1@      @      "@      �?      "@      �?       @               @      �?                      @       @              @      @      @              @      @      �?               @      @       @      @              @       @       @       @      �?              �?       @                      �?               @      $@     `d@      @     �[@      @     �[@      @      ?@               @      @      7@       @      7@      �?       @               @      �?              �?      5@              2@      �?      @      �?      �?      �?                      �?               @      �?                     �S@      �?      �?      �?                      �?      @      J@      @     �H@      @      0@      @      @       @               @      @       @       @              �?       @      �?      �?              �?      �?      �?                      �?               @              (@             �@@       @      @              @       @             �C@      G@      B@      8@      @      ,@      @      �?              �?      @                      *@      >@      $@      <@      @      5@              @      @      @       @      @       @      @                       @      @                      @       @      @       @                      @      @      6@              0@      @      @      @                      @     pq@      b@     �l@     @V@     �j@      Q@               @     �j@     �P@     �H@      C@      E@      C@       @       @      �?              �?       @               @      �?              D@      >@     �@@      <@              @     �@@      7@     �@@      5@      ;@      "@      ;@       @      &@      �?       @      �?              �?       @              "@              0@      @       @      @              @       @              ,@      @      �?      �?              �?      �?              *@       @               @      *@                      �?      @      (@      @      �?              �?      @               @      &@              @       @      @      �?       @      �?                       @      �?      @              @      �?      �?              �?      �?                       @      @       @      @                       @      @             �d@      <@      ;@             @a@      <@     �`@      5@     �`@      ,@     �S@      @      Q@      @     �E@              9@      @      �?       @               @      �?              8@      �?       @      �?              �?       @              0@              &@              K@      &@      K@       @      G@      @      1@      @      ,@      �?       @      �?       @                      �?      (@              @       @      @                       @      =@               @      @      @      @              @      @              @                      @              @      @      @       @              @      @              @      @      @      @      �?              �?      @                       @      1@      5@              "@      1@      (@      @      "@      @       @      @                       @              @      (@      @              �?      (@       @               @      (@              H@      L@      $@      6@      @      �?              �?      @              @      5@              ,@      @      @              @      @      @      @      @      @      �?      @                      �?               @              �?      C@      A@      7@      >@      4@      9@      3@      9@      $@      9@       @      "@      @      @      @      �?      @                      �?              @      @       @      @                       @       @      0@              *@       @      @              @       @              "@              �?              @      @      @                      @      .@      @      ,@      �?      *@              �?      �?      �?                      �?      �?      @              @      �?        r/  tr0  bubhhubh)�r1  }r2  (hhh	h
hNhKhKhG        hh hNhJF<KdhG        hNhG        h<Kh=Kh>h"h#K �r3  h%�r4  Rr5  (KK�r6  hV�C              �?r7  tr8  bhJhZhEC       r9  �r:  Rr;  h^Kh_h`Kh"h#K �r<  h%�r=  Rr>  (KK�r?  hE�C       r@  trA  bK�rB  RrC  }rD  (hKhjMhkh"h#K �rE  h%�rF  RrG  (KM�rH  hr�B88         6                    �?�#i����?�           ��@       #                    a@�zœ���?e            `c@                          �Q@�`�=	�?C            �Y@������������������������       �                     @                          �p@8EGr��?A             Y@                           �?��ɉ�?+            @P@                           �?���J��?!            �I@������������������������       �                     :@	       
       	          ����?`2U0*��?             9@������������������������       �                     4@                           �?z�G�z�?             @������������������������       �                     �?              	          pff�?      �?             @������������������������       �                     �?������������������������       �                     @                           �?@4և���?
             ,@              	             �?$�q-�?	             *@������������������������       �                     (@������������������������       �                     �?������������������������       �                     �?                           �?��R[s�?            �A@                          �d@�����H�?             ;@              	          ����?�nkK�?             7@������������������������       �                     5@              	          pff�?      �?              @������������������������       �                     �?������������������������       �                     �?                          `^@      �?             @������������������������       �                      @������������������������       �                      @       "                    �?      �?              @        !                    �L@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @$       /       	          033�?��
ц��?"             J@%       &                    @H@��Q��?             D@������������������������       �                     @'       *                    �?4���C�?            �@@(       )                   `f@      �?             (@������������������������       �                     "@������������������������       �                     @+       ,                   Pg@���N8�?             5@������������������������       �                     @-       .                    @I@�IєX�?             1@������������������������       �                     �?������������������������       �        
             0@0       5                     P@r�q��?	             (@1       4                    b@�C��2(�?             &@2       3                   `a@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?7       �                    �?�^��[i�?k           �@8       �                    �?h������?�            �r@9       H                    �?���{��?�            @j@:       C       	          @33�?      �?"             H@;       B                    ^@r�q��?             (@<       ?                   0i@�<ݚ�?             "@=       >                   g@      �?              @������������������������       �                     �?������������������������       �                     �?@       A                   `\@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @D       E                   a@������?             B@������������������������       �                     ;@F       G                    `P@�����H�?             "@������������������������       �                      @������������������������       �                     �?I       l       	          ����?$xY+	��?k            @d@J       W                    ]@      �?'             N@K       L                   �Z@���N8�?             5@������������������������       �                     @M       V                   `Z@�����H�?             2@N       S       	          ����?z�G�z�?             $@O       R                    �?      �?              @P       Q                    k@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?T       U                   p`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @X       Y                     D@�99lMt�?            �C@������������������������       �                     @Z       k                   �q@�������?             A@[       h                   �c@r٣����?            �@@\       a                   �h@�>4և��?             <@]       `                   `_@@4և���?	             ,@^       _                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@b       g                    �J@����X�?	             ,@c       f                    �G@�C��2(�?             &@d       e                   �i@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @i       j                    a@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?m       �       	             @��J�x�?D            �Y@n       {                   P`@�7�QJW�?4            �R@o       z       
             �?�&=�w��?&            �J@p       q                    @K@�IєX�?             A@������������������������       �                     0@r       u       	             �?�����H�?             2@s       t                   �U@      �?              @������������������������       �                     �?������������������������       �                     �?v       w                   �^@      �?             0@������������������������       �        	             *@x       y                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     3@|       �       
             �?      �?             6@}       �                    @J@և���X�?	             ,@~       �       	          ����?r�q��?             @       �                   d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �`@      �?              @�       �                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    @H@      �?              @������������������������       �                     @�       �       	             �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     ;@�       �                    �I@�nkK�?9             W@�       �       
             �?�㙢�c�?             7@������������������������       �        
             2@�       �                   �a@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        -            @Q@�       �                    �E@�W��?�            Pq@�       �                   �a@���N8�?#            �O@�       �                   `a@      �?              @������������������������       �                     @������������������������       �                     �?�       �       	             @h㱪��?            �K@������������������������       �                    �J@������������������������       �                      @�       �                    �?�a�4��?�            �j@�       �                   �X@���Q��?d             d@�       �                    �?�C��2(�?             &@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                   pd@
��J���?^            �b@�       �                   P`@xk�2���?N            �_@�       �                   Pa@����X�?(            �Q@�       �                   p@؇���X�?             <@�       �                    �?�nkK�?             7@�       �                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     5@�       �                    @���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   pa@�ՙ/�?             E@������������������������       �                      @�       �                    �?��Q��?             D@�       �                    @L@r�q��?	             (@������������������������       �                     "@�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    _@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    c@և���X�?             <@�       �                    p@���Q��?	             .@�       �                   b@      �?             (@�       �       	          ����?      �?             @�       �                   �i@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    X@�θ�?             *@������������������������       �                     @������������������������       �                     $@�       �                   pi@F�����?&            �L@�       �       	          433�?�X����?             6@������������������������       �        	             *@�       �                   �e@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �       
             �?">�֕�?            �A@�       �                    q@����X�?             @�       �                    �P@r�q��?             @������������������������       �                      @�       �                   �a@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �`@d}h���?             <@�       �                    @�n_Y�K�?
             *@�       �                   �d@���!pc�?	             &@�       �                   �a@�����H�?             "@�       �       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �       	          @33�?��S�ۿ?             .@�       �                   0r@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@�       �                    U@��2(&�?             6@������������������������       �                      @�       �                   �d@P���Q�?             4@�       �                    �?r�q��?             @�       �                     L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        
             ,@�                          hp@����0�?             K@�       �                    �?�+��<��?            �E@������������������������       �                     @�       �                   �O@���Q��?             D@������������������������       �                     $@�       �                   �g@��S���?             >@������������������������       �                     @�       �       
             �?� �	��?             9@�       �                   �`@X�Cc�?             ,@�       �                    [@r�q��?             @������������������������       �                     @�       �                   �k@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    �K@"pc�
�?             &@�       �                   �^@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     &@rI  trJ  bh�h"h#K �rK  h%�rL  RrM  (KMKK�rN  hV�B       `u@     �x@     @]@      C@     @V@      ,@              @     @V@      &@     �O@       @      I@      �?      :@              8@      �?      4@              @      �?      �?              @      �?              �?      @              *@      �?      (@      �?      (@                      �?      �?              :@      "@      8@      @      6@      �?      5@              �?      �?              �?      �?               @       @               @       @               @      @       @       @               @       @                      @      <@      8@      :@      ,@      @              3@      ,@      @      "@              "@      @              0@      @              @      0@      �?              �?      0@               @      $@      �?      $@      �?      @              @      �?                      @      �?              l@      v@      I@     �o@      G@     �d@      @     �F@       @      $@       @      @      �?      �?              �?      �?              �?      @              @      �?                      @      �?     �A@              ;@      �?       @               @      �?             �E@     �]@      >@      >@      @      0@      @               @      0@       @       @      �?      @      �?      @              @      �?                      �?      �?      �?              �?      �?                       @      9@      ,@              @      9@      "@      9@       @      7@      @      *@      �?       @      �?              �?       @              &@              $@      @      $@      �?      @      �?              �?      @              @                      @       @      @       @                      @              �?      *@     @V@      *@      O@       @     �I@       @      @@              0@       @      0@      �?      �?              �?      �?              �?      .@              *@      �?       @      �?                       @              3@      &@      &@       @      @      �?      @      �?      �?              �?      �?                      @      @      �?       @      �?       @                      �?      @              @      @              @      @       @      @                       @              ;@      @      V@      @      3@              2@      @      �?      @                      �?             @Q@     �e@     �Y@      N@      @      @      �?      @                      �?     �J@       @     �J@                       @     �\@     �X@      X@      P@      �?      $@      �?      �?              �?      �?                      "@     �W@      K@      S@     �I@      I@      4@      8@      @      6@      �?      �?      �?              �?      �?              5@               @      @       @                      @      :@      0@               @      :@      ,@      $@       @      "@              �?       @              �?      �?      �?              �?      �?              0@      (@      @      "@      @      "@      @      �?      �?      �?      �?                      �?       @                       @      @              $@      @              @      $@              :@      ?@      .@      @      *@               @      @              @       @              &@      8@      @       @      @      �?       @              @      �?              �?      @                      �?      @      6@      @       @      @       @      �?       @      �?       @      �?                       @              @       @               @              �?      ,@      �?      @      �?                      @              $@      3@      @               @      3@      �?      @      �?      �?      �?      �?                      �?      @              ,@              3@     �A@      3@      8@      @              0@      8@              $@      0@      ,@      @              &@      ,@      "@      @      �?      @              @      �?       @               @      �?               @               @      "@       @       @       @                       @              @              &@rO  trP  bubhhubh)�rQ  }rR  (hhh	h
hNhKhKhG        hh hNhJؽ�hG        hNhG        h<Kh=Kh>h"h#K �rS  h%�rT  RrU  (KK�rV  hV�C              �?rW  trX  bhJhZhEC       rY  �rZ  Rr[  h^Kh_h`Kh"h#K �r\  h%�r]  Rr^  (KK�r_  hE�C       r`  tra  bK�rb  Rrc  }rd  (hKhjM)hkh"h#K �re  h%�rf  Rrg  (KM)�rh  hr�B�@         �                    �?�/�$�y�?�           ��@       U       	          ����?@�0�!��?�            px@       >                    @M@�lg����?Z             `@                           �?     ��?B             X@                          �U@�㙢�c�?             7@������������������������       �                     �?                           �?��2(&�?             6@������������������������       �                     @	                           �?z�G�z�?             .@
                          �`@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?������������������������       �                      @       1                   ``@X~�pX��?5            @R@       ,       
             �? s�n_Y�?$             J@       +                    �?r�q��?             E@       $                    @J@��a�n`�?             ?@              
             �?r�q��?             8@                          @]@r�q��?             @������������������������       �                     @              	             �?�q�q�?             @                           _@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                           �B@r�q��?             2@                          �w@�q�q�?             @������������������������       �                      @������������������������       �                     �?       #                   Pb@��S�ۿ?
             .@               	          ����?      �?             @������������������������       �                      @!       "                   p`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@%       *                   �c@և���X�?             @&       '       
             �?���Q��?             @������������������������       �                     �?(       )                   �g@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     &@-       0                    �?���Q��?             $@.       /       	          @33�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @2       3                   �e@և���X�?             5@������������������������       �                     @4       7                    �?      �?             0@5       6                   �p@�q�q�?             @������������������������       �                     �?������������������������       �                      @8       =                    �?8�Z$���?             *@9       <                   pf@"pc�
�?	             &@:       ;                   8|@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     �?������������������������       �                      @?       T       	          ����?"pc�
�?            �@@@       S                    �?z�G�z�?             >@A       N                    �?�����?             3@B       C       
             �?z�G�z�?             .@������������������������       �                     @D       G                    �?���!pc�?             &@E       F                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?H       M                     P@�<ݚ�?             "@I       L                    �M@      �?              @J       K                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?O       R                    [@      �?             @P       Q                    W@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �        	             &@������������������������       �                     @V       s                    _@���I���?�            `p@W       j                    �?��hJ,�?*             Q@X       ]                    �?ףp=
�?%             N@Y       \                   �]@�<ݚ�?             "@Z       [                    Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @^       i                    @N@�:�]��?            �I@_       f                    @L@������?            �B@`       e                   `]@�FVQ&�?            �@@a       d                    �F@8�Z$���?	             *@b       c                   �X@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �        
             4@g       h                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     ,@k       r       	             @      �?              @l       m                    �?z�G�z�?             @������������������������       �                     �?n       q                   �p@      �?             @o       p                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @t       �                    �R@�'�b�?x            @h@u       �                   �b@     �?w             h@v       {                    �?�(\����?K             ^@w       z                   �r@@4և���?             ,@x       y                   �q@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@|       �                   �z@�O4R���?C            �Z@}       �                    �?�ջ����?A             Z@~                          �c@ ������?*            �O@������������������������       �        &             M@�       �                    �?z�G�z�?             @������������������������       �                      @�       �                   �d@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                    �D@�       �                     L@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�8��8��?,             R@�       �                    `P@�q��/��?            �H@�       �                    �?�C��2(�?             F@�       �                   `o@�X�<ݺ?             B@�       �                   @c@�KM�]�?             3@�       �                    @H@"pc�
�?             &@�       �                   �m@      �?             @������������������������       �                     �?�       �                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     1@�       �                   �_@      �?              @������������������������       �                     @������������������������       �                      @�       �                   �`@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     7@������������������������       �                      @�       �       	             �?0�����?�            pu@�       �                    @L@؇���X�?�            �m@�       �                    �?̫��+�?j             g@�       �                    @<;n,��?c             f@�       �       	          ����?jه��?a            �e@�       �                   `X@ؙ/,T�?\             e@�       �                    ^@����X�?             @������������������������       �                     @������������������������       �                      @�       �                   p@H��%�^�?Z             d@������������������������       �        <            �Z@�       �                    @B@lGts��?            �K@�       �                   Hp@      �?             @������������������������       �                      @������������������������       �                      @�       �                   @g@�:�]��?            �I@�       �                    �? "��u�?             I@�       �                    �? �q�q�?             H@������������������������       �                     >@�       �                    �?�����H�?             2@������������������������       �                     "@�       �                   pa@�<ݚ�?             "@������������������������       �                     @�       �                   �q@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �H@z�G�z�?             @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �d@      �?              @������������������������       �                     @�       �       
             �?���Q��?             @�       �                    �G@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �       	          ��������0�?"             K@������������������������       �                     @�       �                   �O@�\�u��?!            �I@�       �                    �?���|���?             &@�       �                    �?����X�?             @������������������������       �                     �?�       �                    `@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     �?�       �                     P@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �M@R���Q�?             D@�       �       
             �?X�<ݚ�?             "@�       �                    @z�G�z�?             @�       �                    �L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    �?      �?             @�       �                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                   �W@��� ��?             ?@������������������������       �                     �?�       �                   �c@ףp=
�?             >@�       �                    �?@4և���?             <@������������������������       �                     (@�       �                    b@      �?
             0@������������������������       �                     &@�       �                   @h@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?�                          �?&RN���?G            @Z@�       �                   `X@�q�q�?             8@������������������������       �                      @�       �                    �L@��2(&�?             6@�       �                    �?      �?             0@������������������������       �                     @�       �                   �b@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?�                          �?�q�q�?             @�                          `c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                        �c@2lK����?6            @T@            	          pff�?����>4�?%             L@                        �_@X�Cc�?             <@      	                  �Q@@�0�!��?
             1@            	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @
                         @M@@4և���?             ,@������������������������       �                      @                         @N@r�q��?             @������������������������       �                     �?������������������������       �                     @                        0q@���|���?	             &@                         @M@      �?              @                         �?      �?             @������������������������       �                     �?������������������������       �                     @                        (p@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                         �?h�����?             <@                         �N@���N8�?             5@������������������������       �        	             0@                        �`@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @      &      	             @`�Q��?             9@       #                   �?�S����?             3@!      "                   �L@��S�ۿ?	             .@������������������������       �                     ,@������������������������       �                     �?$      %                  �d@      �?             @������������������������       �                      @������������������������       �                      @'      (      	          ���
@r�q��?             @������������������������       �                     @������������������������       �                     �?ri  trj  bh�h"h#K �rk  h%�rl  Rrm  (KM)KK�rn  hV�B�        t@     �y@     @Q@      t@      H@     @T@      E@      K@      3@      @              �?      3@      @      @              (@      @      (@      �?      (@                      �?               @      7@      I@      &@     �D@      @     �A@      @      8@      @      4@      �?      @              @      �?       @      �?      �?      �?                      �?              �?      @      .@       @      �?       @                      �?      �?      ,@      �?      @               @      �?      �?              �?      �?                      &@      @      @      @       @      �?               @       @       @                       @               @              &@      @      @      @      �?      @                      �?              @      (@      "@              @      (@      @      �?       @      �?                       @      &@       @      "@       @      "@      �?      "@                      �?              �?       @              @      ;@      @      8@      @      *@      @      (@              @      @       @      �?      �?              �?      �?               @      @      �?      @      �?       @               @      �?                      @      �?              @      �?      �?      �?      �?                      �?       @                      &@              @      5@      n@      $@      M@      @      K@       @      @       @      �?              �?       @                      @      @     �G@      @     �@@       @      ?@       @      &@       @      �?              �?       @                      $@              4@       @       @       @                       @              ,@      @      @      �?      @              �?      �?      @      �?      �?      �?                      �?               @      @              &@     �f@      "@     �f@      @     @]@      �?      *@      �?      @              @      �?                      "@       @      Z@      �?     �Y@      �?      O@              M@      �?      @               @      �?       @      �?                       @             �D@      �?      �?              �?      �?              @     �P@      @     �E@      @      D@       @      A@       @      1@       @      "@       @       @      �?              �?       @               @      �?                      @               @              1@       @      @              @       @               @      @              @       @                      7@       @             `o@      W@     �i@      A@      e@      .@     `d@      *@      d@      (@     �c@      &@       @      @              @       @             `c@      @     �Z@             �H@      @       @       @               @       @             �G@      @     �G@      @      G@       @      >@              0@       @      "@              @       @      @              �?       @      �?                       @      �?      �?              �?      �?                      �?      @      �?       @               @      �?      �?              �?      �?      �?                      �?       @      �?       @                      �?      @       @      @              @       @       @       @               @       @              �?             �A@      3@              @     �A@      0@      @      @       @      @      �?              �?      @              @      �?               @       @              �?       @      �?              �?       @              ?@      "@      @      @      �?      @      �?       @               @      �?                       @      @      �?       @      �?              �?       @              �?              ;@      @              �?      ;@      @      :@       @      (@              ,@       @      &@              @       @      @                       @      �?      �?              �?      �?             �G@      M@      3@      @               @      3@      @      .@      �?      @              (@      �?      (@                      �?      @       @      �?       @      �?                       @      @              <@     �J@      &@     �F@      $@      2@      @      ,@       @      �?              �?       @              �?      *@               @      �?      @      �?                      @      @      @      @      @      �?      @      �?                      @      @      �?      @                      �?      @              �?      ;@      �?      4@              0@      �?      @      �?                      @              @      1@       @      0@      @      ,@      �?      ,@                      �?       @       @       @                       @      �?      @              @      �?        ro  trp  bubhhubh)�rq  }rr  (hhh	h
hNhKhKhG        hh hNhJX��vhG        hNhG        h<Kh=Kh>h"h#K �rs  h%�rt  Rru  (KK�rv  hV�C              �?rw  trx  bhJhZhEC       ry  �rz  Rr{  h^Kh_h`Kh"h#K �r|  h%�r}  Rr~  (KK�r  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjK�hkh"h#K �r�  h%�r�  Rr�  (KK�r�  hr�B2         x       	          ����?���
%�?�           ��@                          �O@���u�J�?�            �v@                           �?�S����?&            �L@                          �Z@��R[s�?            �A@������������������������       �                      @                          @[@�q�q�?             ;@������������������������       �                      @              
             �? �o_��?             9@	       
                    �?@�0�!��?	             1@������������������������       �                     &@                          �a@      �?             @                          �]@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                           �?      �?              @                          �]@      �?             @������������������������       �                      @������������������������       �                      @                          �\@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     6@       3                   �`@�d�����?�             s@       &                    �?B� ��?)            �Q@                           �?�I�w�"�?             C@                          0i@�����H�?             "@������������������������       �                     �?������������������������       �                      @                          �Y@�c�Α�?             =@������������������������       �                      @        !                   �Y@�<ݚ�?             ;@������������������������       �                     @"       #                    �?      �?             8@������������������������       �                     �?$       %       	          ����?���}<S�?
             7@������������������������       �                     5@������������������������       �                      @'       2                    �?     ��?             @@(       +                   �X@d}h���?             <@)       *                   @\@      �?             @������������������������       �                     @������������������������       �                     @,       -                    �?��2(&�?             6@������������������������       �                     @.       /                   `c@z�G�z�?             .@������������������������       �                     &@0       1                   pn@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @4       ?                    �?�?�m�?�            @m@5       <                   �d@������?5            �T@6       7                   �`@pY���D�?3            �S@������������������������       �        )             P@8       ;                   @o@�r����?
             .@9       :                   �n@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @=       >                    q@�q�q�?             @������������������������       �                      @������������������������       �                     �?@       S                    �?�|�ʒ�?c             c@A       H                    �?X�<ݚ�?            �F@B       G       	             �?r�q��?
             2@C       D                    @F@z�G�z�?             .@������������������������       �                     @E       F                   f@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @I       P                    �?��}*_��?             ;@J       M                   �c@��H�}�?             9@K       L                   �a@@4և���?             ,@������������������������       �                     *@������������������������       �                     �?N       O                    t@���!pc�?             &@������������������������       �                      @������������������������       �                     @Q       R                    �?      �?              @������������������������       �                     �?������������������������       �                     �?T       o       	            �?$	4�}�?H            �Z@U       n                   �d@Hm_!'1�?A            �X@V       g                    �L@      �??             X@W       X                   0n@Pq�����?5            @U@������������������������       �                    �F@Y       f                    �?ףp=
�?             D@Z       [                    �?$�q-�?            �C@������������������������       �                     =@\       ]                   �n@�z�G��?             $@������������������������       �                      @^       _       
             �?      �?              @������������������������       �                     �?`       e                    f@؇���X�?             @a       b                    \@�q�q�?             @������������������������       �                     �?c       d                   @p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?h       m                   hr@"pc�
�?
             &@i       j       
             �?ףp=
�?	             $@������������������������       �                     @k       l                   0a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @p       w                   xp@X�<ݚ�?             "@q       r                   �`@�q�q�?             @������������������������       �                     @s       v                    �?�q�q�?             @t       u       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @y       �                    �?|��T+[�?�            Pw@z       �                    �?ؓ!'�s�?�            `n@{       �                   @]@"pc�
�?             F@|       }                    �?z�G�z�?             @������������������������       �                      @~              	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �J@��-�=��?            �C@�       �                    �?�	j*D�?             *@�       �       	          ����?      �?              @������������������������       �                      @�       �       	          ����?�q�q�?             @������������������������       �                      @�       �                   h@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     :@�       �       
             �?������?�            �h@�       �                    �?�U�e?Ƕ?d            �b@�       �                    �H@      �?             @@������������������������       �                     �?�       �       	             @�g�y��?             ?@������������������������       �                     8@�       �       	          ���@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                   �Q@Xc!J�ƴ?M            �]@������������������������       �                     �?�       �                    `R@ȑ����?L            @]@�       �                   �U@ �^�@̩?K             ]@������������������������       �                     �?�       �                    q@�]���?J            �\@�       �                    I@�q�q�??             X@�       �                   P`@�g�y��?             ?@������������������������       �                     :@�       �                    @M@z�G�z�?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        (            @P@�       �                   8q@�}�+r��?             3@�       �                   @b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             1@������������������������       �                     �?�       �       	          ����?Hm_!'1�?$            �H@�       �       	          033�?��s����?             5@�       �                    @H@�����H�?	             "@������������������������       �                     �?������������������������       �                      @�       �                    �N@      �?             (@������������������������       �                      @�       �                   �`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     <@�       �                    �?
j*D>�?L            @`@�       �                    �?XB���?             =@������������������������       �                     (@�       �                   �g@�IєX�?             1@�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             .@�       �                    �F@zP1�?:            @Y@�       �                    �?�<ݚ�?             "@������������������������       �                      @�       �       	              @����X�?             @������������������������       �                     @������������������������       �                      @�       �                   �b@��<b���?5             W@�       �                   P`@��IF�E�?#            �P@�       �                    �?�t����?             1@�       �                   �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �K@d}h���?             ,@������������������������       �                     $@�       �                   @a@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   pb@@9G��?            �H@������������������������       �                     @@�       �                    �?�t����?             1@������������������������       �                     "@�       �                   �a@      �?              @�       �                    �M@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    b@      �?             :@�       �                    �?\X��t�?             7@�       �       
             �?؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                    d@      �?             0@�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �h@�C��2(�?             &@�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hV�BP       0s@     �z@      m@      `@      "@      H@      "@      :@               @      "@      2@       @              @      2@      @      ,@              &@      @      @      @      �?              �?      @                       @      @      @       @       @       @                       @       @       @               @       @                      6@      l@      T@      ?@     �C@      "@      =@      �?       @      �?                       @       @      5@       @              @      5@      @              @      5@      �?               @      5@              5@       @              6@      $@      6@      @      @      @      @                      @      3@      @      @              (@      @      &@              �?      @      �?                      @              @      h@     �D@     �S@      @     @S@       @      P@              *@       @      @       @      @                       @       @              �?       @               @      �?             �\@     �B@      4@      9@      @      .@      @      (@              @      @      @              @      @                      @      1@      $@      0@      "@      *@      �?      *@                      �?      @       @               @      @              �?      �?      �?                      �?     �W@      (@     �V@       @     �V@      @     @T@      @     �F@              B@      @      B@      @      =@              @      @               @      @      �?      �?              @      �?       @      �?      �?              �?      �?      �?                      �?      @                      �?      "@       @      "@      �?      @               @      �?       @                      �?              �?               @      @      @       @      @              @       @      �?      �?      �?      �?                      �?      �?              @             �R@     �r@      3@      l@       @      B@      @      �?       @               @      �?              �?       @              @     �A@      @      "@      @      @       @               @      @               @       @       @       @                       @              @              :@      &@     �g@      @     �a@       @      >@      �?              �?      >@              8@      �?      @      �?                      @      @     @\@      �?              @     @\@      @     @\@      �?               @     @\@      �?     �W@      �?      >@              :@      �?      @              @      �?      �?      �?                      �?             @P@      �?      2@      �?      �?      �?                      �?              1@      �?              @     �F@      @      1@      �?       @      �?                       @      @      "@               @      @      �?      @                      �?              <@     �K@     �R@      <@      �?      (@              0@      �?      �?      �?      �?                      �?      .@              ;@     �R@      @       @       @              @       @      @                       @      4@      R@      @     �M@      @      (@       @      �?              �?       @              @      &@              $@      @      �?              �?      @               @     �G@              @@       @      .@              "@       @      @       @      �?              �?       @                      @      *@      *@      $@      *@      @      �?              �?      @              @      (@      @       @               @      @              �?      $@      �?       @               @      �?                       @      @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ���EhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjMhkh"h#K �r�  h%�r�  Rr�  (KM�r�  hr�B9         �       	          033�?�r,��?�           ��@       u                    �?H;N	�	�?�             x@                          @E@��;�\`�?�             u@                           Z@�99lMt�?            �C@������������������������       �                     @                          �\@�������?             A@������������������������       �        
             2@       	                     I@     ��?             0@������������������������       �                     @
                           �?      �?
             (@������������������������       �                     �?                           �P@"pc�
�?	             &@������������������������       �                      @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @       Z                   pq@�$�����?�            �r@       /                   `_@��A���?�             n@       *                   �^@���Q��?            �F@                          �k@�����?             C@                          �\@�㙢�c�?             7@              
             �?���Q��?             @������������������������       �                     @������������������������       �                      @                          0a@�X�<ݺ?             2@������������������������       �                     &@                           �?؇���X�?             @������������������������       �                      @                          �f@z�G�z�?             @������������������������       �                     �?������������������������       �                     @        )                    b@��S���?             .@!       "                    �?���|���?             &@������������������������       �                     @#       (                   @`@�q�q�?             @$       %       
             �?z�G�z�?             @������������������������       �                     �?&       '                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @+       .                    j@؇���X�?             @,       -                    _@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @0       G                    �?��-�=��?y            `h@1       4                    �?�BbΊ�?!             M@2       3                   �n@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?5       6                   �[@p�v>��?            �G@������������������������       �                     @7       >                   �b@d}h���?             E@8       9                   Pj@�����H�?             ;@������������������������       �                     3@:       =                   pk@      �?              @;       <                   0a@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @?       @                    @E@���Q��?
             .@������������������������       �                     �?A       B       
             �?X�Cc�?	             ,@������������������������       �                     @C       F                    �?      �?             $@D       E       	             �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @H       Q       	          pff�?���Z�?X             a@I       J       
             �?��v$���?N            �^@������������������������       �        A             Y@K       L                    �?�C��2(�?             6@������������������������       �                      @M       N                    j@؇���X�?             ,@������������������������       �                      @O       P                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     @R       S                   �_@z�G�z�?
             .@������������������������       �                     @T       Y                   0m@      �?              @U       X       
             �?���Q��?             @V       W                   c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @[       h                   s@���b���?"            �L@\       _       
             �?     ��?             @@]       ^       	          @33�?�����H�?             "@������������������������       �                      @������������������������       �                     �?`       c                    �C@
;&����?             7@a       b                    r@؇���X�?             @������������������������       �                     @������������������������       �                     �?d       e                    @E@     ��?	             0@������������������������       �                     @f       g                    �?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @i       j                    �@@�J�4�?             9@������������������������       �                     �?k       l                    �?      �?             8@������������������������       �        	             0@m       t                   8|@      �?              @n       s                   �d@����X�?             @o       p                    �H@�q�q�?             @������������������������       �                     �?q       r                    �M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?v       �                    �?Fx$(�?#             I@w       x                    �?��S�ۿ?             >@������������������������       �                     @y       z                   ``@�>����?             ;@������������������������       �        
             .@{       �       	          833�?r�q��?             (@|              	          ����?�<ݚ�?             "@}       ~                   �p@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �W@R���Q�?             4@������������������������       �                     �?�       �                   �U@�KM�]�?             3@������������������������       �                     �?�       �                    �?�X�<ݺ?             2@�       �                   �m@r�q��?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@�       �                   �b@д>��C�?�            �u@�       �                   P`@܍�l�p�?�             r@�       �                    �?�P��G7�?Q            @]@�       �                    �?JyK���??            �U@�       �       	          pff�?�n_Y�K�?             *@�       �                     K@X�<ݚ�?             "@�       �                   �_@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    V@x!'ǯ�?8            �R@������������������������       �                     �?�       �       
             �?��W��?7            @R@�       �                   Hs@X�;�^o�?*            �K@�       �                    �E@`�H�/��?'            �I@������������������������       �                      @�       �                   @^@X�EQ]N�?"            �E@�       �                   �Y@д>��C�?             =@������������������������       �                     @�       �                   �j@z�G�z�?             9@�       �       	             �?�eP*L��?
             &@������������������������       �                     �?�       �       	          `ff�?���Q��?	             $@�       �       
             �?z�G�z�?             @������������������������       �                     �?�       �                   �^@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?���Q��?             @������������������������       �                      @�       �                    @L@�q�q�?             @������������������������       �                     �?�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             ,@������������������������       �                     ,@�       �       	          @33�?      �?             @������������������������       �                      @������������������������       �                      @�       �       	          033�?b�2�tk�?             2@�       �       	          033�?�<ݚ�?             "@�       �                   �[@����X�?             @�       �                   �Y@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    n@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �       	             �?X�<ݚ�?             "@������������������������       �                     @�       �       	             @�q�q�?             @�       �                     D@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   @`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     >@�       �                    @Pt�nٔ�?e            �e@�       �                   �b@��AV���?b            �d@�       �                   �a@�L��ȕ?4            @W@������������������������       �        .            �T@�       �                     K@�C��2(�?             &@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �       
             �?,N�_� �?.            �R@�       �                    �?�h����?!             L@�       �                    `@�?�|�?            �B@������������������������       �                     7@�       �                    �H@@4և���?             ,@�       �                    �G@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     3@�       �                   �u@�<ݚ�?             2@�       �                   P`@@�0�!��?             1@������������������������       �        	             &@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   0c@      �?&             M@������������������������       �                      @�       �                    �G@���H.�?"             I@�       �                    @B@z�G�z�?
             .@������������������������       �                     �?�       �                    V@؇���X�?	             ,@������������������������       �                      @������������������������       �                     (@�       �                   �e@��R[s�?            �A@�       �                     L@���Q��?             @������������������������       �                     �?�       �                    �O@      �?             @������������������������       �                     @������������������������       �                     �?�       �       	          ����?z�G�z�?             >@������������������������       �                      @�                         �d@���!pc�?             6@�             	          033�?ҳ�wY;�?             1@�                           �?�q�q�?             @�       �                    �?�q�q�?             @�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                        �m@"pc�
�?             &@������������������������       �                      @������������������������       �                     "@������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMKK�r�  hV�BP       �t@     Py@     �p@     @]@     @o@     �U@      ,@      9@      @              "@      9@              2@      "@      @              @      "@      @              �?      "@       @       @              �?       @      �?                       @     �m@     �N@     @i@      C@      ;@      2@      :@      (@      3@      @       @      @              @       @              1@      �?      &@              @      �?       @              @      �?              �?      @              @       @      @      @      @               @      @      �?      @              �?      �?      @              @      �?              �?                      @      �?      @      �?      �?      �?                      �?              @     �e@      4@     �E@      .@      $@      �?      $@                      �?     �@@      ,@              @     �@@      "@      8@      @      3@              @      @      �?      @              @      �?              @              "@      @              �?      "@      @      @              @      @      @      @              @      @               @             �`@      @      ^@       @      Y@              4@       @       @              (@       @       @              @       @               @      @              (@      @      @              @      @       @      @       @      �?              �?       @                       @      @              A@      7@      *@      3@      �?       @               @      �?              (@      &@      �?      @              @      �?              &@      @      @              @      @      @                      @      5@      @              �?      5@      @      0@              @      @      @       @      �?       @              �?      �?      �?      �?                      �?      @                      �?      3@      ?@       @      <@              @       @      9@              .@       @      $@       @      @      �?      @              @      �?              �?                      @      1@      @              �?      1@       @              �?      1@      �?      @      �?      @               @      �?      �?              �?      �?      �?                      �?      (@              N@      r@      ?@     0p@      7@     �W@      7@      P@       @      @      @      @      �?      @      �?                      @      @              @              .@     �M@      �?              ,@     �M@      @      H@      @      G@               @      @      C@      @      8@              @      @      4@      @      @      �?              @      @      �?      @              �?      �?      @              @      �?              @       @       @              �?       @              �?      �?      �?              �?      �?                      ,@              ,@       @       @       @                       @      @      &@       @      @       @      @      �?      �?              �?      �?              �?      @      �?                      @               @      @      @      @               @      @      �?      @      �?                      @      �?      �?              �?      �?                      >@       @     �d@      @      d@      �?      W@             �T@      �?      $@      �?      �?      �?                      �?              "@      @     @Q@      �?     �K@      �?      B@              7@      �?      *@      �?      @              @      �?                      @              3@      @      ,@      @      ,@              &@      @      @      @                      @      �?               @      @       @                      @      =@      =@       @              5@      =@      (@      @              �?      (@       @               @      (@              "@      :@      @       @              �?      @      �?      @                      �?      @      8@               @      @      0@      @      &@      @       @      �?       @      �?      �?      �?                      �?              �?      @               @      "@       @                      "@              @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ:9)bhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjK�hkh"h#K �r�  h%�r�  Rr�  (KK�r�  hr�Bh3         8                    �?T8���?�           ��@       -                    �?�<ݚ��?_             b@                          `a@���B���?V            @`@                           �?`Jj��?=            @W@                           �D@     ��?             @@������������������������       �                     �?                           �?��� ��?             ?@������������������������       �                     @	                          �`@�J�4�?             9@
              	          ����?      �?             8@������������������������       �        	             ,@                          �[@�z�G��?             $@              	          `ff�?      �?              @������������������������       �                     �?������������������������       �                     �?                           �I@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     �?                           �?��v$���?)            �N@������������������������       �        !             H@                           �?$�q-�?             *@������������������������       �                     @                          p@r�q��?             @������������������������       �                     @������������������������       �                     �?       $                   �b@��+��?            �B@                           �?����X�?             5@������������������������       �                     &@       #                    @���Q��?             $@       "                   �a@և���X�?             @        !                    �N@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @%       ,       	          ���@      �?             0@&       '                    �?$�q-�?	             *@������������������������       �                      @(       )                    �?z�G�z�?             @������������������������       �                     @*       +                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @.       7                   �s@և���X�?	             ,@/       6                   `b@���!pc�?             &@0       5       	          `ff�?      �?              @1       2                    @I@����X�?             @������������������������       �                     �?3       4                     @r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @9       �                    �?2� J��?p           p�@:       �       	          033�?��׸���?            }@;       \                   `_@�w��#��?�            @o@<       =                    Z@b�2�tk�?-             R@������������������������       �                     @>       O                   `c@ҳ�wY;�?*             Q@?       H                    �?     ��?             @@@       G                     Q@�J�4�?             9@A       F                    �?      �?             8@B       C                   �_@@�0�!��?             1@������������������������       �                     @D       E                    `@�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?I       N       	             �?����X�?             @J       M                   @_@r�q��?             @K       L                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?P       W                   �[@      �?             B@Q       V                    `@�LQ�1	�?             7@R       S                    k@�n_Y�K�?             *@������������������������       �                     @T       U                    �N@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     $@X       [                    �K@�θ�?	             *@Y       Z                    �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @]       ~                   �o@dWp,��?k            @f@^       m                   Pi@�HP��a�?B            @[@_       `                   �\@�GN�z�?             F@������������������������       �                      @a       l                    �?�X�<ݺ?             B@b       c                    @I@�<ݚ�?             "@������������������������       �                     @d       e                     K@�q�q�?             @������������������������       �                     �?f       g                   @`@z�G�z�?             @������������������������       �                      @h       i                     M@�q�q�?             @������������������������       �                     �?j       k                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ;@n       o       
             �?$�q-�?(            @P@������������������������       �                     "@p       }       
             �?4և����?!             L@q       |                    @ףp=
�?             I@r       {                   �f@Hm_!'1�?            �H@s       v                   �a@`�q�0ܴ?            �G@t       u                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @w       x       	            �?��Y��]�?            �D@������������������������       �                    �C@y       z                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @       �                   h}@bKv���?)            @Q@�       �                    @K@҄��?(            �P@�       �       	          ����?l��
I��?!             K@�       �                    �?"Ae���?            �G@�       �                   �t@      �?
             (@�       �                    @I@ףp=
�?             $@������������������������       �                      @�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �       
             �?z�G�z�?            �A@�       �                    f@��� ��?             ?@�       �                    �? 	��p�?             =@�       �                   @p@���}<S�?             7@������������������������       �                      @������������������������       �                     5@������������������������       �                     @������������������������       �                      @�       �                     E@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �c@�q�q�?             (@�       �                   �`@X�<ݚ�?             "@������������������������       �                     @�       �                     L@z�G�z�?             @�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                     F@�e/
�?�             k@�       �                   �b@П[;U��?             =@�       �                   �l@@4և���?
             ,@������������������������       �                     $@�       �                   �n@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     .@�       �                   `j@a��_�?p            `g@�       �                   0`@Xny��?&            �N@������������������������       �                    �B@�       �                   p`@�q�q�?             8@������������������������       �                     @�       �                    �?��s����?             5@�       �       	          ����?      �?             0@������������������������       �                     @�       �                    �G@�q�q�?             (@������������������������       �                     �?�       �                   @_@���!pc�?             &@�       �                   �W@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?�Ń��̧?J            �_@�       �                   0a@p���?9             Y@������������������������       �                    �F@�       �                    @K@h㱪��?            �K@�       �                    �?�KM�]�?             3@�       �                     J@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?�IєX�?
             1@�       �                   �m@      �?             @������������������������       �                      @�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@������������������������       �                     B@�       �                    �H@ ��WV�?             :@�       �                   �l@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     3@�       �                    _@�z�6�?V             _@�       �       	          `ff@(;L]n�?+             N@������������������������       �        )            �L@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �P@      �?+             P@�       �                   �c@`��}3��?$            �J@�       �       	          433�?"pc�
�?             F@�       �                     M@�z�G��?             $@������������������������       �                     @������������������������       �                     @�       �                    y@г�wY;�?             A@������������������������       �                     @@�       �                     L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                   �p@���|���?             &@�       �                   pm@؇���X�?             @������������������������       �                     @�       �                   �^@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   c@      �?             @������������������������       �                      @�       �                   @e@      �?              @������������������������       �                     �?������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hV�B�       �t@     @y@     @\@      ?@     @Z@      9@     �U@      @      ;@      @              �?      ;@      @      @              5@      @      5@      @      ,@              @      @      �?      �?              �?      �?              @       @               @      @                      �?      N@      �?      H@              (@      �?      @              @      �?      @                      �?      2@      3@      @      .@              &@      @      @      @      @      �?      @              @      �?               @              @              (@      @      (@      �?       @              @      �?      @              �?      �?              �?      �?                      @       @      @       @      @      @      @      @       @              �?      @      �?      @                      �?              �?      @                      @      k@     Pw@     �g@     0q@     �d@     @U@      <@      F@      @              8@      F@      @      :@      @      5@      @      5@      @      ,@              @      @      @      @                      @              @      �?               @      @      �?      @      �?      @              @      �?                       @      �?              2@      2@      .@       @      @       @              @      @      @              @      @              $@              @      $@      @      @              @      @                      @      a@     �D@     �W@      .@      A@      $@               @      A@       @      @       @      @              @       @              �?      @      �?       @               @      �?      �?              �?      �?      �?                      �?      ;@              N@      @      "@             �I@      @     �F@      @     �F@      @     �F@       @      @      �?              �?      @              D@      �?     �C@              �?      �?      �?                      �?               @              �?      @             �E@      :@     �E@      7@      C@      0@      ?@      0@      @      "@      �?      "@               @      �?      �?              �?      �?               @              <@      @      ;@      @      ;@       @      5@       @               @      5@              @                       @      �?      @      �?                      @      @              @      @      @      @      @              �?      @      �?      �?              �?      �?                      @              @              @      :@     �g@      0@      *@      �?      *@              $@      �?      @      �?                      @      .@              $@      f@      @      K@             �B@      @      1@      @              @      1@      @      (@              @      @       @      �?              @       @       @      �?       @                      �?      �?      @      �?                      @              @      @     �^@       @     �X@             �F@       @     �J@       @      1@      �?      �?              �?      �?              �?      0@      �?      @               @      �?      �?              �?      �?                      *@              B@      �?      9@      �?      @              @      �?                      3@      :@     �X@       @      M@             �L@       @      �?              �?       @              8@      D@      1@      B@       @      B@      @      @      @                      @      �?     �@@              @@      �?      �?              �?      �?              "@              @      @      @      �?      @              @      �?              �?      @              �?      @               @      �?      �?      �?                      �?r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�BHzhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjMhkh"h#K �r�  h%�r�  Rr�  (KM�r�  hr�B88         �       	          ����?�[��N�?�           ��@                           �?��)��?�            �v@                           _@*
;&���?5             W@                           �J@�n_Y�K�?             *@                           [@      �?             @������������������������       �                     �?������������������������       �                     @                           `R@�<ݚ�?             "@	       
                    @      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?                          @d@l{��b��?-            �S@                          �Q@@-�_ .�?*            �R@������������������������       �                     �?                           �?���(-�?)            @R@              
             �?r�q��?             (@������������������������       �                     $@������������������������       �                      @                           �?��v$���?!            �N@������������������������       �                    �J@                          �`@      �?              @������������������������       �                     @                          @q@      �?              @������������������������       �                     �?������������������������       �                     �?                           f@���Q��?             @������������������������       �                      @������������������������       �                     @       Q                    �?N{�T6�?�            0q@       .                   `_@3k���?E            @\@        '                   �j@�q��/��?             G@!       "                   �Z@�˹�m��?             C@������������������������       �                     .@#       $                     E@�LQ�1	�?             7@������������������������       �                      @%       &                   �Z@���N8�?             5@������������������������       �                     �?������������������������       �                     4@(       -       	             �?      �?              @)       ,                    �?؇���X�?             @*       +                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?/       F                   ``@�2�,��?(            �P@0       1                    �?�q�q�?             E@������������������������       �                     "@2       3                   �V@4���C�?            �@@������������������������       �                      @4       =                   �b@� �	��?             9@5       <                   �x@d}h���?             ,@6       ;                   �a@8�Z$���?             *@7       :                   pk@����X�?             @8       9                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?>       ?                    �B@���!pc�?             &@������������������������       �                      @@       A                     E@�����H�?             "@������������������������       �                     @B       E                   �]@z�G�z�?             @C       D                    @F@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?G       P       	          pff�?z�G�z�?             9@H       K                    �?�LQ�1	�?             7@I       J                   �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?L       M                   �n@P���Q�?
             4@������������������������       �                     0@N       O                    d@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @R       e                   `_@ʰ-M���?a            @d@S       d                    �?����e��?            �@@T       a       
             �?�q�q�?             >@U       X                    �?�+e�X�?             9@V       W                   `V@      �?             @������������������������       �                     �?������������������������       �                     @Y       `                   @_@؇���X�?             5@Z       _                    �L@�z�G��?             $@[       \                    �?      �?              @������������������������       �                     @]       ^                    @G@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@b       c                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @f       �                   �g@(L���?M             `@g       �                    @ ��P0�?L            �_@h       k                   @[@�=|+g��?E            @\@i       j       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @l       u                    @L@,�+�C�?C            �[@m       r       	            �?X;��?7            @V@n       q                    �A@ qP��B�?5            �U@o       p                   Pb@"pc�
�?             &@������������������������       �                      @������������������������       �                     "@������������������������       �        -            �R@s       t                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?v                          Ps@���N8�?             5@w       z                    `@z�G�z�?             4@x       y                   Pk@���Q��?             @������������������������       �                      @������������������������       �                     @{       ~                   �`@��S�ۿ?	             .@|       }                    `@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@������������������������       �                     �?�       �                    �M@և���X�?             ,@������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                    �?ByL5���?�            �v@�       �                    �?���>4��?(             L@�       �                    �?�<ݚ�?             B@�       �                   �_@r�q��?             >@�       �                    �P@�q�q�?             "@�       �       	             �?      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                   �a@�����?             5@�       �                    �?؇���X�?
             ,@�       �                   h@      �?              @������������������������       �                     �?�       �                    a@؇���X�?             @������������������������       �                     @�       �       	          033@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                     L@      �?             @������������������������       �                     @������������������������       �                     @�       �       	          ����?ףp=
�?             4@�       �                   �g@      �?              @������������������������       �                     �?�       �                   �Z@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@�       �                    �E@���?�            ps@�       �       	          ����?�	j*D�?             :@�       �                   xt@     ��?             0@�       �                    �?�r����?             .@������������������������       �        
             *@������������������������       �                      @������������������������       �                     �?�       �                    @C@      �?             $@������������������������       �                     @�       �                    h@����X�?             @������������������������       �                      @������������������������       �                     @�       �                   �v@4z:V��?�            �q@�       �                    _@xzY���?�            �q@�       �                   ``@(;L]n�?Z            �b@�       �                    �?�>����?!             K@������������������������       �                     C@�       �       	             @      �?	             0@�       �                   �]@؇���X�?             ,@�       �                   @_@$�q-�?             *@������������������������       �                      @�       �                   �X@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?�q�q�?9             X@�       �                   �c@$�q-�?             *@������������������������       �                     $@�       �                   �d@�q�q�?             @�       �                    `@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �        2            �T@�       �                    �?�����D�?R            @`@�       �                   Pi@��8��)�?;            �W@�       �       
             �?d}h���?             <@�       �                    a@��2(&�?             6@�       �                   i@      �?             (@�       �                    �?ףp=
�?             $@������������������������       �                     @�       �                   P`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@�       �       	          033�?      �?             @������������������������       �                     @������������������������       �                     @�       �                    �?���7�?+            �P@�       �                   �c@�]0��<�?&            �N@�       �                   �[@ _�@�Y�?#             M@�       �                    �I@r�q��?             @�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     J@�       �                   �d@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                      @�       �                    c@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	          ����?�q�q�?             B@�       �                   �k@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                   �b@������?             ;@�       �                    �?�t����?             1@�       �                    @��S�ۿ?
             .@������������������������       �                     $@�       �                   �k@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    b@      �?             $@�       �       
             �?����X�?             @�       �                    �K@r�q��?             @�       �                   Pm@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   ``@���Q��?             @������������������������       �                      @�                           �J@�q�q�?             @������������������������       �                     �?������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMKK�r�  hV�B       �s@     Pz@      o@     �]@     �S@      ,@      @       @      @      �?              �?      @               @      @      �?      @              @      �?              �?             @R@      @     �Q@      @              �?     �Q@      @      $@       @      $@                       @      N@      �?     �J@              @      �?      @              �?      �?              �?      �?              @       @               @      @             @e@     @Z@     �C@     �R@      @     �D@      @     �A@              .@      @      4@       @              �?      4@      �?                      4@       @      @      �?      @      �?      �?              �?      �?                      @      �?              A@     �@@      ,@      <@              "@      ,@      3@               @      ,@      &@      &@      @      &@       @      @       @      �?       @               @      �?              @              @                      �?      @       @       @              �?       @              @      �?      @      �?      @      �?                      @              �?      4@      @      4@      @      �?       @               @      �?              3@      �?      0@              @      �?              �?      @                       @     ``@      ?@      4@      *@      4@      $@      3@      @      �?      @      �?                      @      2@      @      @      @      @      �?      @              @      �?      @                      �?               @      &@              �?      @      �?                      @              @     �[@      2@     �[@      0@     �Y@      $@      �?       @      �?                       @     �Y@       @     �U@      @      U@       @      "@       @               @      "@             �R@               @      �?       @                      �?      0@      @      0@      @       @      @       @                      @      ,@      �?      �?      �?      �?                      �?      *@                      �?       @      @              @       @                       @     @P@     �r@      :@      >@       @      <@      @      9@      @      @       @      @       @                      @      �?               @      3@       @      (@       @      @      �?              �?      @              @      �?      �?      �?                      �?              @              @      @      @      @                      @      2@       @      @       @              �?      @      �?              �?      @              (@             �C@      q@       @      2@      @      *@       @      *@              *@       @              �?              @      @              @      @       @               @      @              ?@     �o@      =@     `o@      @      b@      @      I@              C@      @      (@       @      (@      �?      (@               @      �?      @      �?                      @      �?               @              �?     �W@      �?      (@              $@      �?       @      �?      �?      �?                      �?              �?             �T@      8@     �Z@      "@     @U@      @      6@      @      3@      @      "@      �?      "@              @      �?      @              @      �?               @                      $@      @      @              @      @              @     �O@       @     �M@      �?     �L@      �?      @      �?       @      �?                       @              @              J@      �?       @      �?                       @      �?      @               @      �?       @               @      �?              .@      5@       @      �?              �?       @              @      4@       @      .@      �?      ,@              $@      �?      @      �?                      @      �?      �?              �?      �?              @      @       @      @      �?      @      �?       @      �?                       @              @      �?              @               @      @               @       @      �?              �?       @        r�  tr�  bubhhubehhub.